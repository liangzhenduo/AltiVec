//===============================================================================
//  File Name       : AltiVecUnit.v
//  File Revision   : 1.0
//  Date            : 2015/3/30
//  Author          : wangjie
//  Email           : ycyquick@foxmail.com
//  ----------------------------------------------------------------------------
//  Description     : Vector Registers (for students)
//  Function        : three read ports, no need latency five write ports, 1 latency
//  ----------------------------------------------------------------------------
// Copyright (c) 2015,Tianjin University.
//               No.92 Weijin Road , Nankai District, Tianjin, 300072, China
// Tianjin University Confidential Proprietary
//===============================================================================

module RegisterFile(
                 clk,
                 rst_n,
                 in_AReadRegisterEnable,
                 in_AReadRegister,
                 in_BReadRegisterEnable,
                 in_BReadRegister,
                 in_CReadRegisterEnable,
                 in_CReadRegister,
                 in_ZeroWriteRegister,
                 in_ZeroWriteData,
                 in_ZeroWriteRegisterEnable,
                 in_FirstWriteRegisterEnable,
                 in_FirstWriteRegister,
                 in_FirstWriteData,
                 in_SecondWriteRegisterEnable,
                 in_SecondWriteRegister,
                 in_SecondWriteData,
                 in_ThirdWriteRegisterEnable,
                 in_ThirdWriteRegister,
                 in_ThirdWriteData,
                 in_FourthWriteRegisterEnable,
                 in_FourthWriteRegister,
                 in_FourthWriteData,
                 in_FifthWriteRegisterEnable,
                 in_FifthWriteRegister,
                 in_FifthWriteData,

                 out_AReadData,
                 out_BReadData,
                 out_CReadData
                 );

//===============================================================================
//input and output declaration
//===============================================================================
input            clk;
input            rst_n;
//3 read port
//first read port
input            in_AReadRegisterEnable;
input    [0:  4] in_AReadRegister;
//second read port
input            in_BReadRegisterEnable;
input    [0:  4] in_BReadRegister;
//third read port
input            in_CReadRegisterEnable;
input    [0:  4] in_CReadRegister;

//Load/Store write port
input    [0: 15] in_ZeroWriteRegisterEnable;
input    [0:  4] in_ZeroWriteRegister;
input    [0:127] in_ZeroWriteData;
//PU write port
input            in_FirstWriteRegisterEnable;
input    [0:  4] in_FirstWriteRegister;
input    [0:127] in_FirstWriteData;
//VSFX write port
input            in_SecondWriteRegisterEnable;
input    [0:  4] in_SecondWriteRegister;
input    [0:127] in_SecondWriteData;
//VCFX write port
input            in_ThirdWriteRegisterEnable;
input    [0:  4] in_ThirdWriteRegister;
input    [0:127] in_ThirdWriteData;
//VFPU write port
input            in_FourthWriteRegisterEnable;
input    [0:  4] in_FourthWriteRegister;
input    [0:127] in_FourthWriteData;
//VSCR write port
input            in_FifthWriteRegisterEnable;
input    [0:  4] in_FifthWriteRegister;
input    [0: 31] in_FifthWriteData;

//first read data out
output   [0:127] out_AReadData;
//second read data out
output   [0:127] out_BReadData;
//third read data out
output   [0:127] out_CReadData;

//---------------------------------------------------------------------
//Internal signals declaration
//-----------------------------------------------------------------------
// | ------------   write reg0 mask   ------------ |
// | bit0       | bit1 | bit2 | bit  | bit4 | bit5 |
// | Load/Store | PU   | VSFX | VCFX | VFPU | VSCR |
wire     [0:  5] Reg0WriteMask;
wire     [0:  5] Reg1WriteMask;
wire     [0:  5] Reg2WriteMask;
wire     [0:  5] Reg3WriteMask;
wire     [0:  5] Reg4WriteMask;
wire     [0:  5] Reg5WriteMask;
wire     [0:  5] Reg6WriteMask;
wire     [0:  5] Reg7WriteMask;
wire     [0:  5] Reg8WriteMask;
wire     [0:  5] Reg9WriteMask;
wire     [0:  5] Reg10WriteMask;
wire     [0:  5] Reg11WriteMask;
wire     [0:  5] Reg12WriteMask;
wire     [0:  5] Reg13WriteMask;
wire     [0:  5] Reg14WriteMask;
wire     [0:  5] Reg15WriteMask;
wire     [0:  5] Reg16WriteMask;
wire     [0:  5] Reg17WriteMask;
wire     [0:  5] Reg18WriteMask;
wire     [0:  5] Reg19WriteMask;
wire     [0:  5] Reg20WriteMask;
wire     [0:  5] Reg21WriteMask;
wire     [0:  5] Reg22WriteMask;
wire     [0:  5] Reg23WriteMask;
wire     [0:  5] Reg24WriteMask;
wire     [0:  5] Reg25WriteMask;
wire     [0:  5] Reg26WriteMask;
wire     [0:  5] Reg27WriteMask;
wire     [0:  5] Reg28WriteMask;
wire     [0:  5] Reg29WriteMask;
wire     [0:  5] Reg30WriteMask;
wire     [0:  5] Reg31WriteMask;

//===============================================================================
//internal registers
//===============================================================================
//reg style declaration of output signal
reg      [0:127] out_AReadData;
reg      [0:127] out_BReadData;
reg      [0:127] out_CReadData;
reg      [0:127] Reg0;
reg      [0:127] Reg1;
reg      [0:127] Reg2;
reg      [0:127] Reg3;
reg      [0:127] Reg4;
reg      [0:127] Reg5;
reg      [0:127] Reg6;
reg      [0:127] Reg7;
reg      [0:127] Reg8;
reg      [0:127] Reg9;
reg      [0:127] Reg10;
reg      [0:127] Reg11;
reg      [0:127] Reg12;
reg      [0:127] Reg13;
reg      [0:127] Reg14;
reg      [0:127] Reg15;
reg      [0:127] Reg16;
reg      [0:127] Reg17;
reg      [0:127] Reg18;
reg      [0:127] Reg19;
reg      [0:127] Reg20;
reg      [0:127] Reg21;
reg      [0:127] Reg22;
reg      [0:127] Reg23;
reg      [0:127] Reg24;
reg      [0:127] Reg25;
reg      [0:127] Reg26;
reg      [0:127] Reg27;
reg      [0:127] Reg28;
reg      [0:127] Reg29;
reg      [0:127] Reg30;
reg      [0:127] Reg31;

//===============================================================================
//write  registers
//===============================================================================
//generate write mask signal
assign Reg0WriteMask  = {{(|in_ZeroWriteRegisterEnable) && ( in_ZeroWriteRegister   == 5'd0  )},
                         { in_FirstWriteRegisterEnable  && ( in_FirstWriteRegister  == 5'd0  )},
                         { in_SecondWriteRegisterEnable && ( in_SecondWriteRegister == 5'd0  )},
                         { in_ThirdWriteRegisterEnable  && ( in_ThirdWriteRegister  == 5'd0  )},
                         { in_FourthWriteRegisterEnable && ( in_FourthWriteRegister == 5'd0  )},
                         { in_FifthWriteRegisterEnable  && ( in_FifthWriteRegister  == 5'd0  )}};
assign Reg1WriteMask  = {{(|in_ZeroWriteRegisterEnable) && ( in_ZeroWriteRegister   == 5'd1  )},
                         { in_FirstWriteRegisterEnable  && ( in_FirstWriteRegister  == 5'd1  )},
                         { in_SecondWriteRegisterEnable && ( in_SecondWriteRegister == 5'd1  )},
                         { in_ThirdWriteRegisterEnable  && ( in_ThirdWriteRegister  == 5'd1  )},
                         { in_FourthWriteRegisterEnable && ( in_FourthWriteRegister == 5'd1  )},
                         { in_FifthWriteRegisterEnable  && ( in_FifthWriteRegister  == 5'd1  )}};
assign Reg2WriteMask  = {{(|in_ZeroWriteRegisterEnable) && ( in_ZeroWriteRegister   == 5'd2  )},
                         { in_FirstWriteRegisterEnable  && ( in_FirstWriteRegister  == 5'd2  )},
                         { in_SecondWriteRegisterEnable && ( in_SecondWriteRegister == 5'd2  )},
                         { in_ThirdWriteRegisterEnable  && ( in_ThirdWriteRegister  == 5'd2  )},
                         { in_FourthWriteRegisterEnable && ( in_FourthWriteRegister == 5'd2  )},
                         { in_FifthWriteRegisterEnable  && ( in_FifthWriteRegister  == 5'd2  )}};
assign Reg3WriteMask  = {{(|in_ZeroWriteRegisterEnable) && ( in_ZeroWriteRegister   == 5'd3  )},
                         { in_FirstWriteRegisterEnable  && ( in_FirstWriteRegister  == 5'd3  )},
                         { in_SecondWriteRegisterEnable && ( in_SecondWriteRegister == 5'd3  )},
                         { in_ThirdWriteRegisterEnable  && ( in_ThirdWriteRegister  == 5'd3  )},
                         { in_FourthWriteRegisterEnable && ( in_FourthWriteRegister == 5'd3  )},
                         { in_FifthWriteRegisterEnable  && ( in_FifthWriteRegister  == 5'd3  )}};
assign Reg4WriteMask  = {{(|in_ZeroWriteRegisterEnable) && ( in_ZeroWriteRegister   == 5'd4  )},
                         { in_FirstWriteRegisterEnable  && ( in_FirstWriteRegister  == 5'd4  )},
                         { in_SecondWriteRegisterEnable && ( in_SecondWriteRegister == 5'd4  )},
                         { in_ThirdWriteRegisterEnable  && ( in_ThirdWriteRegister  == 5'd4  )},
                         { in_FourthWriteRegisterEnable && ( in_FourthWriteRegister == 5'd4  )},
                         { in_FifthWriteRegisterEnable  && ( in_FifthWriteRegister  == 5'd4  )}};
assign Reg5WriteMask  = {{(|in_ZeroWriteRegisterEnable) && ( in_ZeroWriteRegister   == 5'd5  )},
                         { in_FirstWriteRegisterEnable  && ( in_FirstWriteRegister  == 5'd5  )},
                         { in_SecondWriteRegisterEnable && ( in_SecondWriteRegister == 5'd5  )},
                         { in_ThirdWriteRegisterEnable  && ( in_ThirdWriteRegister  == 5'd5  )},
                         { in_FourthWriteRegisterEnable && ( in_FourthWriteRegister == 5'd5  )},
                         { in_FifthWriteRegisterEnable  && ( in_FifthWriteRegister  == 5'd5  )}};
assign Reg6WriteMask  = {{(|in_ZeroWriteRegisterEnable) && ( in_ZeroWriteRegister   == 5'd6  )},
                         { in_FirstWriteRegisterEnable  && ( in_FirstWriteRegister  == 5'd6  )},
                         { in_SecondWriteRegisterEnable && ( in_SecondWriteRegister == 5'd6  )},
                         { in_ThirdWriteRegisterEnable  && ( in_ThirdWriteRegister  == 5'd6  )},
                         { in_FourthWriteRegisterEnable && ( in_FourthWriteRegister == 5'd6  )},
                         { in_FifthWriteRegisterEnable  && ( in_FifthWriteRegister  == 5'd6  )}};
assign Reg7WriteMask  = {{(|in_ZeroWriteRegisterEnable) && ( in_ZeroWriteRegister   == 5'd7  )},
                         { in_FirstWriteRegisterEnable  && ( in_FirstWriteRegister  == 5'd7  )},
                         { in_SecondWriteRegisterEnable && ( in_SecondWriteRegister == 5'd7  )},
                         { in_ThirdWriteRegisterEnable  && ( in_ThirdWriteRegister  == 5'd7  )},
                         { in_FourthWriteRegisterEnable && ( in_FourthWriteRegister == 5'd7  )},
                         { in_FifthWriteRegisterEnable  && ( in_FifthWriteRegister  == 5'd7  )}};
assign Reg8WriteMask  = {{(|in_ZeroWriteRegisterEnable) && ( in_ZeroWriteRegister   == 5'd8  )},
                         { in_FirstWriteRegisterEnable  && ( in_FirstWriteRegister  == 5'd8  )},
                         { in_SecondWriteRegisterEnable && ( in_SecondWriteRegister == 5'd8  )},
                         { in_ThirdWriteRegisterEnable  && ( in_ThirdWriteRegister  == 5'd8  )},
                         { in_FourthWriteRegisterEnable && ( in_FourthWriteRegister == 5'd8  )},
                         { in_FifthWriteRegisterEnable  && ( in_FifthWriteRegister  == 5'd8  )}};
assign Reg9WriteMask  = {{(|in_ZeroWriteRegisterEnable) && ( in_ZeroWriteRegister   == 5'd9  )},
                         { in_FirstWriteRegisterEnable  && ( in_FirstWriteRegister  == 5'd9  )},
                         { in_SecondWriteRegisterEnable && ( in_SecondWriteRegister == 5'd9  )},
                         { in_ThirdWriteRegisterEnable  && ( in_ThirdWriteRegister  == 5'd9  )},
                         { in_FourthWriteRegisterEnable && ( in_FourthWriteRegister == 5'd9  )},
                         { in_FifthWriteRegisterEnable  && ( in_FifthWriteRegister  == 5'd9  )}};
assign Reg10WriteMask = {{(|in_ZeroWriteRegisterEnable) && ( in_ZeroWriteRegister   == 5'd10 )},
                         { in_FirstWriteRegisterEnable  && ( in_FirstWriteRegister  == 5'd10 )},
                         { in_SecondWriteRegisterEnable && ( in_SecondWriteRegister == 5'd10 )},
                         { in_ThirdWriteRegisterEnable  && ( in_ThirdWriteRegister  == 5'd10 )},
                         { in_FourthWriteRegisterEnable && ( in_FourthWriteRegister == 5'd10 )},
                         { in_FifthWriteRegisterEnable  && ( in_FifthWriteRegister  == 5'd10 )}};
assign Reg11WriteMask = {{(|in_ZeroWriteRegisterEnable) && ( in_ZeroWriteRegister   == 5'd11 )},
                         { in_FirstWriteRegisterEnable  && ( in_FirstWriteRegister  == 5'd11 )},
                         { in_SecondWriteRegisterEnable && ( in_SecondWriteRegister == 5'd11 )},
                         { in_ThirdWriteRegisterEnable  && ( in_ThirdWriteRegister  == 5'd11 )},
                         { in_FourthWriteRegisterEnable && ( in_FourthWriteRegister == 5'd11 )},
                         { in_FifthWriteRegisterEnable  && ( in_FifthWriteRegister  == 5'd11 )}};
assign Reg12WriteMask = {{(|in_ZeroWriteRegisterEnable) && ( in_ZeroWriteRegister   == 5'd12 )},
                         { in_FirstWriteRegisterEnable  && ( in_FirstWriteRegister  == 5'd12 )},
                         { in_SecondWriteRegisterEnable && ( in_SecondWriteRegister == 5'd12 )},
                         { in_ThirdWriteRegisterEnable  && ( in_ThirdWriteRegister  == 5'd12 )},
                         { in_FourthWriteRegisterEnable && ( in_FourthWriteRegister == 5'd12 )},
                         { in_FifthWriteRegisterEnable  && ( in_FifthWriteRegister  == 5'd12 )}};
assign Reg13WriteMask = {{(|in_ZeroWriteRegisterEnable) && ( in_ZeroWriteRegister   == 5'd13 )},
                         { in_FirstWriteRegisterEnable  && ( in_FirstWriteRegister  == 5'd13 )},
                         { in_SecondWriteRegisterEnable && ( in_SecondWriteRegister == 5'd13 )},
                         { in_ThirdWriteRegisterEnable  && ( in_ThirdWriteRegister  == 5'd13 )},
                         { in_FourthWriteRegisterEnable && ( in_FourthWriteRegister == 5'd13 )},
                         { in_FifthWriteRegisterEnable  && ( in_FifthWriteRegister  == 5'd13 )}};
assign Reg14WriteMask = {{(|in_ZeroWriteRegisterEnable) && ( in_ZeroWriteRegister   == 5'd14 )},
                         { in_FirstWriteRegisterEnable  && ( in_FirstWriteRegister  == 5'd14 )},
                         { in_SecondWriteRegisterEnable && ( in_SecondWriteRegister == 5'd14 )},
                         { in_ThirdWriteRegisterEnable  && ( in_ThirdWriteRegister  == 5'd14 )},
                         { in_FourthWriteRegisterEnable && ( in_FourthWriteRegister == 5'd14 )},
                         { in_FifthWriteRegisterEnable  && ( in_FifthWriteRegister  == 5'd14 )}};
assign Reg15WriteMask = {{(|in_ZeroWriteRegisterEnable) && ( in_ZeroWriteRegister   == 5'd15 )},
                         { in_FirstWriteRegisterEnable  && ( in_FirstWriteRegister  == 5'd15 )},
                         { in_SecondWriteRegisterEnable && ( in_SecondWriteRegister == 5'd15 )},
                         { in_ThirdWriteRegisterEnable  && ( in_ThirdWriteRegister  == 5'd15 )},
                         { in_FourthWriteRegisterEnable && ( in_FourthWriteRegister == 5'd15 )},
                         { in_FifthWriteRegisterEnable  && ( in_FifthWriteRegister  == 5'd15 )}};
assign Reg16WriteMask = {{(|in_ZeroWriteRegisterEnable) && ( in_ZeroWriteRegister   == 5'd16 )},
                         { in_FirstWriteRegisterEnable  && ( in_FirstWriteRegister  == 5'd16 )},
                         { in_SecondWriteRegisterEnable && ( in_SecondWriteRegister == 5'd16 )},
                         { in_ThirdWriteRegisterEnable  && ( in_ThirdWriteRegister  == 5'd16 )},
                         { in_FourthWriteRegisterEnable && ( in_FourthWriteRegister == 5'd16 )},
                         { in_FifthWriteRegisterEnable  && ( in_FifthWriteRegister  == 5'd16 )}};
assign Reg17WriteMask = {{(|in_ZeroWriteRegisterEnable) && ( in_ZeroWriteRegister   == 5'd17 )},
                         { in_FirstWriteRegisterEnable  && ( in_FirstWriteRegister  == 5'd17 )},
                         { in_SecondWriteRegisterEnable && ( in_SecondWriteRegister == 5'd17 )},
                         { in_ThirdWriteRegisterEnable  && ( in_ThirdWriteRegister  == 5'd17 )},
                         { in_FourthWriteRegisterEnable && ( in_FourthWriteRegister == 5'd17 )},
                         { in_FifthWriteRegisterEnable  && ( in_FifthWriteRegister  == 5'd17 )}};
assign Reg18WriteMask = {{(|in_ZeroWriteRegisterEnable) && ( in_ZeroWriteRegister   == 5'd18 )},
                         { in_FirstWriteRegisterEnable  && ( in_FirstWriteRegister  == 5'd18 )},
                         { in_SecondWriteRegisterEnable && ( in_SecondWriteRegister == 5'd18 )},
                         { in_ThirdWriteRegisterEnable  && ( in_ThirdWriteRegister  == 5'd18 )},
                         { in_FourthWriteRegisterEnable && ( in_FourthWriteRegister == 5'd18 )},
                         { in_FifthWriteRegisterEnable  && ( in_FifthWriteRegister  == 5'd18 )}};
assign Reg19WriteMask = {{(|in_ZeroWriteRegisterEnable) && ( in_ZeroWriteRegister   == 5'd19 )},
                         { in_FirstWriteRegisterEnable  && ( in_FirstWriteRegister  == 5'd19 )},
                         { in_SecondWriteRegisterEnable && ( in_SecondWriteRegister == 5'd19 )},
                         { in_ThirdWriteRegisterEnable  && ( in_ThirdWriteRegister  == 5'd19 )},
                         { in_FourthWriteRegisterEnable && ( in_FourthWriteRegister == 5'd19 )},
                         { in_FifthWriteRegisterEnable  && ( in_FifthWriteRegister  == 5'd19 )}};
assign Reg20WriteMask = {{(|in_ZeroWriteRegisterEnable) && ( in_ZeroWriteRegister   == 5'd20 )},
                         { in_FirstWriteRegisterEnable  && ( in_FirstWriteRegister  == 5'd20 )},
                         { in_SecondWriteRegisterEnable && ( in_SecondWriteRegister == 5'd20 )},
                         { in_ThirdWriteRegisterEnable  && ( in_ThirdWriteRegister  == 5'd20 )},
                         { in_FourthWriteRegisterEnable && ( in_FourthWriteRegister == 5'd20 )},
                         { in_FifthWriteRegisterEnable  && ( in_FifthWriteRegister  == 5'd20 )}};
assign Reg21WriteMask = {{(|in_ZeroWriteRegisterEnable) && ( in_ZeroWriteRegister   == 5'd21 )},
                         { in_FirstWriteRegisterEnable  && ( in_FirstWriteRegister  == 5'd21 )},
                         { in_SecondWriteRegisterEnable && ( in_SecondWriteRegister == 5'd21 )},
                         { in_ThirdWriteRegisterEnable  && ( in_ThirdWriteRegister  == 5'd21 )},
                         { in_FourthWriteRegisterEnable && ( in_FourthWriteRegister == 5'd21 )},
                         { in_FifthWriteRegisterEnable  && ( in_FifthWriteRegister  == 5'd21 )}};
assign Reg22WriteMask = {{(|in_ZeroWriteRegisterEnable) && ( in_ZeroWriteRegister   == 5'd22 )},
                         { in_FirstWriteRegisterEnable  && ( in_FirstWriteRegister  == 5'd22 )},
                         { in_SecondWriteRegisterEnable && ( in_SecondWriteRegister == 5'd22 )},
                         { in_ThirdWriteRegisterEnable  && ( in_ThirdWriteRegister  == 5'd22 )},
                         { in_FourthWriteRegisterEnable && ( in_FourthWriteRegister == 5'd22 )},
                         { in_FifthWriteRegisterEnable  && ( in_FifthWriteRegister  == 5'd22 )}};
assign Reg23WriteMask = {{(|in_ZeroWriteRegisterEnable) && ( in_ZeroWriteRegister   == 5'd23 )},
                         { in_FirstWriteRegisterEnable  && ( in_FirstWriteRegister  == 5'd23 )},
                         { in_SecondWriteRegisterEnable && ( in_SecondWriteRegister == 5'd23 )},
                         { in_ThirdWriteRegisterEnable  && ( in_ThirdWriteRegister  == 5'd23 )},
                         { in_FourthWriteRegisterEnable && ( in_FourthWriteRegister == 5'd23 )},
                         { in_FifthWriteRegisterEnable  && ( in_FifthWriteRegister  == 5'd23 )}};
assign Reg24WriteMask = {{(|in_ZeroWriteRegisterEnable) && ( in_ZeroWriteRegister   == 5'd24 )},
                         { in_FirstWriteRegisterEnable  && ( in_FirstWriteRegister  == 5'd24 )},
                         { in_SecondWriteRegisterEnable && ( in_SecondWriteRegister == 5'd24 )},
                         { in_ThirdWriteRegisterEnable  && ( in_ThirdWriteRegister  == 5'd24 )},
                         { in_FourthWriteRegisterEnable && ( in_FourthWriteRegister == 5'd24 )},
                         { in_FifthWriteRegisterEnable  && ( in_FifthWriteRegister  == 5'd24 )}};
assign Reg25WriteMask = {{(|in_ZeroWriteRegisterEnable) && ( in_ZeroWriteRegister   == 5'd25 )},
                         { in_FirstWriteRegisterEnable  && ( in_FirstWriteRegister  == 5'd25 )},
                         { in_SecondWriteRegisterEnable && ( in_SecondWriteRegister == 5'd25 )},
                         { in_ThirdWriteRegisterEnable  && ( in_ThirdWriteRegister  == 5'd25 )},
                         { in_FourthWriteRegisterEnable && ( in_FourthWriteRegister == 5'd25 )},
                         { in_FifthWriteRegisterEnable  && ( in_FifthWriteRegister  == 5'd25 )}};
assign Reg26WriteMask = {{(|in_ZeroWriteRegisterEnable) && ( in_ZeroWriteRegister   == 5'd26 )},
                         { in_FirstWriteRegisterEnable  && ( in_FirstWriteRegister  == 5'd26 )},
                         { in_SecondWriteRegisterEnable && ( in_SecondWriteRegister == 5'd26 )},
                         { in_ThirdWriteRegisterEnable  && ( in_ThirdWriteRegister  == 5'd26 )},
                         { in_FourthWriteRegisterEnable && ( in_FourthWriteRegister == 5'd26 )},
                         { in_FifthWriteRegisterEnable  && ( in_FifthWriteRegister  == 5'd26 )}};
assign Reg27WriteMask = {{(|in_ZeroWriteRegisterEnable) && ( in_ZeroWriteRegister   == 5'd27 )},
                         { in_FirstWriteRegisterEnable  && ( in_FirstWriteRegister  == 5'd27 )},
                         { in_SecondWriteRegisterEnable && ( in_SecondWriteRegister == 5'd27 )},
                         { in_ThirdWriteRegisterEnable  && ( in_ThirdWriteRegister  == 5'd27 )},
                         { in_FourthWriteRegisterEnable && ( in_FourthWriteRegister == 5'd27 )},
                         { in_FifthWriteRegisterEnable  && ( in_FifthWriteRegister  == 5'd27 )}};
assign Reg28WriteMask = {{(|in_ZeroWriteRegisterEnable) && ( in_ZeroWriteRegister   == 5'd28 )},
                         { in_FirstWriteRegisterEnable  && ( in_FirstWriteRegister  == 5'd28 )},
                         { in_SecondWriteRegisterEnable && ( in_SecondWriteRegister == 5'd28 )},
                         { in_ThirdWriteRegisterEnable  && ( in_ThirdWriteRegister  == 5'd28 )},
                         { in_FourthWriteRegisterEnable && ( in_FourthWriteRegister == 5'd28 )},
                         { in_FifthWriteRegisterEnable  && ( in_FifthWriteRegister  == 5'd28 )}};
assign Reg29WriteMask = {{(|in_ZeroWriteRegisterEnable) && ( in_ZeroWriteRegister   == 5'd29 )},
                         { in_FirstWriteRegisterEnable  && ( in_FirstWriteRegister  == 5'd29 )},
                         { in_SecondWriteRegisterEnable && ( in_SecondWriteRegister == 5'd29 )},
                         { in_ThirdWriteRegisterEnable  && ( in_ThirdWriteRegister  == 5'd29 )},
                         { in_FourthWriteRegisterEnable && ( in_FourthWriteRegister == 5'd29 )},
                         { in_FifthWriteRegisterEnable  && ( in_FifthWriteRegister  == 5'd29)}};
assign Reg30WriteMask = {{(|in_ZeroWriteRegisterEnable) && ( in_ZeroWriteRegister   == 5'd30 )},
                         { in_FirstWriteRegisterEnable  && ( in_FirstWriteRegister  == 5'd30 )},
                         { in_SecondWriteRegisterEnable && ( in_SecondWriteRegister == 5'd30 )},
                         { in_ThirdWriteRegisterEnable  && ( in_ThirdWriteRegister  == 5'd30 )},
                         { in_FourthWriteRegisterEnable && ( in_FourthWriteRegister == 5'd30 )},
                         { in_FifthWriteRegisterEnable  && ( in_FifthWriteRegister  == 5'd30 )}};
assign Reg31WriteMask = {{(|in_ZeroWriteRegisterEnable) && ( in_ZeroWriteRegister   == 5'd31 )},
                         { in_FirstWriteRegisterEnable  && ( in_FirstWriteRegister  == 5'd31 )},
                         { in_SecondWriteRegisterEnable && ( in_SecondWriteRegister == 5'd31 )},
                         { in_ThirdWriteRegisterEnable  && ( in_ThirdWriteRegister  == 5'd31 )},
                         { in_FourthWriteRegisterEnable && ( in_FourthWriteRegister == 5'd31 )},
                         { in_FifthWriteRegisterEnable  && ( in_FifthWriteRegister  == 5'd31 )}};

//===============================================================================
//read  A registers
//===============================================================================
always @ ( Reg0  or Reg1  or Reg2  or Reg3  or Reg4  or Reg5  or Reg6  or Reg7  or
           Reg8  or Reg9  or Reg10 or Reg11 or Reg12 or Reg13 or Reg14 or Reg15 or
           Reg16 or Reg17 or Reg18 or Reg19 or Reg20 or Reg21 or Reg22 or Reg23 or
           Reg24 or Reg25 or Reg26 or Reg27 or Reg28 or Reg29 or Reg30 or Reg31 or
           in_AReadRegisterEnable or in_AReadRegister )
  if(in_AReadRegisterEnable)
  begin
    case(in_AReadRegister)
      5'd0    : out_AReadData = Reg0;
      5'd1    : out_AReadData = Reg1;
      5'd2    : out_AReadData = Reg2;
      5'd3    : out_AReadData = Reg3;
      5'd4    : out_AReadData = Reg4;
      5'd5    : out_AReadData = Reg5;
      5'd6    : out_AReadData = Reg6;
      5'd7    : out_AReadData = Reg7;
      5'd8    : out_AReadData = Reg8;
      5'd9    : out_AReadData = Reg9;
      5'd10   : out_AReadData = Reg10;
      5'd11   : out_AReadData = Reg11;
      5'd12   : out_AReadData = Reg12;
      5'd13   : out_AReadData = Reg13;
      5'd14   : out_AReadData = Reg14;
      5'd15   : out_AReadData = Reg15;
      5'd16   : out_AReadData = Reg16;
      5'd17   : out_AReadData = Reg17;
      5'd18   : out_AReadData = Reg18;
      5'd19   : out_AReadData = Reg19;
      5'd20   : out_AReadData = Reg20;
      5'd21   : out_AReadData = Reg21;
      5'd22   : out_AReadData = Reg22;
      5'd23   : out_AReadData = Reg23;
      5'd24   : out_AReadData = Reg24;
      5'd25   : out_AReadData = Reg25;
      5'd26   : out_AReadData = Reg26;
      5'd27   : out_AReadData = Reg27;
      5'd28   : out_AReadData = Reg28;
      5'd29   : out_AReadData = Reg29;
      5'd30   : out_AReadData = Reg30;
      default : out_AReadData = Reg31;
    endcase
  end
  else
    out_AReadData = 128'b0;

//===============================================================================
//read  B registers
//===============================================================================
always @ ( Reg0  or Reg1  or Reg2  or Reg3  or Reg4  or Reg5  or Reg6  or Reg7  or
           Reg8  or Reg9  or Reg10 or Reg11 or Reg12 or Reg13 or Reg14 or Reg15 or
           Reg16 or Reg17 or Reg18 or Reg19 or Reg20 or Reg21 or Reg22 or Reg23 or
           Reg24 or Reg25 or Reg26 or Reg27 or Reg28 or Reg29 or Reg30 or Reg31 or
           in_BReadRegisterEnable or in_BReadRegister )
  if(in_BReadRegisterEnable)
  begin
    case(in_BReadRegister)
      5'd0    : out_BReadData = Reg0;
      5'd1    : out_BReadData = Reg1;
      5'd2    : out_BReadData = Reg2;
      5'd3    : out_BReadData = Reg3;
      5'd4    : out_BReadData = Reg4;
      5'd5    : out_BReadData = Reg5;
      5'd6    : out_BReadData = Reg6;
      5'd7    : out_BReadData = Reg7;
      5'd8    : out_BReadData = Reg8;
      5'd9    : out_BReadData = Reg9;
      5'd10   : out_BReadData = Reg10;
      5'd11   : out_BReadData = Reg11;
      5'd12   : out_BReadData = Reg12;
      5'd13   : out_BReadData = Reg13;
      5'd14   : out_BReadData = Reg14;
      5'd15   : out_BReadData = Reg15;
      5'd16   : out_BReadData = Reg16;
      5'd17   : out_BReadData = Reg17;
      5'd18   : out_BReadData = Reg18;
      5'd19   : out_BReadData = Reg19;
      5'd20   : out_BReadData = Reg20;
      5'd21   : out_BReadData = Reg21;
      5'd22   : out_BReadData = Reg22;
      5'd23   : out_BReadData = Reg23;
      5'd24   : out_BReadData = Reg24;
      5'd25   : out_BReadData = Reg25;
      5'd26   : out_BReadData = Reg26;
      5'd27   : out_BReadData = Reg27;
      5'd28   : out_BReadData = Reg28;
      5'd29   : out_BReadData = Reg29;
      5'd30   : out_BReadData = Reg30;
      default : out_BReadData = Reg31;
    endcase
  end
  else
    out_BReadData = 128'b0;

//===============================================================================
//read  C registers
//===============================================================================
always @ ( Reg0  or Reg1  or Reg2  or Reg3  or Reg4  or Reg5  or Reg6  or Reg7  or
           Reg8  or Reg9  or Reg10 or Reg11 or Reg12 or Reg13 or Reg14 or Reg15 or
           Reg16 or Reg17 or Reg18 or Reg19 or Reg20 or Reg21 or Reg22 or Reg23 or
           Reg24 or Reg25 or Reg26 or Reg27 or Reg28 or Reg29 or Reg30 or Reg31 or
           in_CReadRegisterEnable or in_CReadRegister )
  if(in_CReadRegisterEnable)
  begin
    case(in_CReadRegister)
      5'd0    : out_CReadData = Reg0;
      5'd1    : out_CReadData = Reg1;
      5'd2    : out_CReadData = Reg2;
      5'd3    : out_CReadData = Reg3;
      5'd4    : out_CReadData = Reg4;
      5'd5    : out_CReadData = Reg5;
      5'd6    : out_CReadData = Reg6;
      5'd7    : out_CReadData = Reg7;
      5'd8    : out_CReadData = Reg8;
      5'd9    : out_CReadData = Reg9;
      5'd10   : out_CReadData = Reg10;
      5'd11   : out_CReadData = Reg11;
      5'd12   : out_CReadData = Reg12;
      5'd13   : out_CReadData = Reg13;
      5'd14   : out_CReadData = Reg14;
      5'd15   : out_CReadData = Reg15;
      5'd16   : out_CReadData = Reg16;
      5'd17   : out_CReadData = Reg17;
      5'd18   : out_CReadData = Reg18;
      5'd19   : out_CReadData = Reg19;
      5'd20   : out_CReadData = Reg20;
      5'd21   : out_CReadData = Reg21;
      5'd22   : out_CReadData = Reg22;
      5'd23   : out_CReadData = Reg23;
      5'd24   : out_CReadData = Reg24;
      5'd25   : out_CReadData = Reg25;
      5'd26   : out_CReadData = Reg26;
      5'd27   : out_CReadData = Reg27;
      5'd28   : out_CReadData = Reg28;
      5'd29   : out_CReadData = Reg29;
      5'd30   : out_CReadData = Reg30;
      default : out_CReadData = Reg31;
    endcase
  end
  else
    out_CReadData = 128'b0;

//write data to registerfile according to write mask signal
//0  1  2    3    4    5
//LS PU VSFX VCFX VFPU VALU

//write Reg0
always @ ( posedge clk or negedge rst_n )
begin
  if( !rst_n )
  begin
    Reg0 <= 128'h0;
  end
  else if ( | Reg0WriteMask )
  begin
    case ( Reg0WriteMask )
      6'b100000 : begin
					if (in_ZeroWriteRegisterEnable[0])
						Reg0[  0:  7] <= in_ZeroWriteData[  0:  7];
					if (in_ZeroWriteRegisterEnable[1])
						Reg0[  8: 15] <= in_ZeroWriteData[  8: 15];
					if (in_ZeroWriteRegisterEnable[2])
						Reg0[ 16: 23] <= in_ZeroWriteData[ 16: 23];
					if (in_ZeroWriteRegisterEnable[3])
						Reg0[ 24: 31] <= in_ZeroWriteData[ 24: 31];
					if (in_ZeroWriteRegisterEnable[4])
						Reg0[ 32: 39] <= in_ZeroWriteData[ 32: 39];
					if (in_ZeroWriteRegisterEnable[5])
						Reg0[ 40: 47] <= in_ZeroWriteData[ 40: 47];
					if (in_ZeroWriteRegisterEnable[6])
						Reg0[ 48: 55] <= in_ZeroWriteData[ 48: 55];
					if (in_ZeroWriteRegisterEnable[7])
						Reg0[ 56: 63] <= in_ZeroWriteData[ 56: 63];
					if (in_ZeroWriteRegisterEnable[8])
						Reg0[ 64: 71] <= in_ZeroWriteData[ 64: 71];
					if (in_ZeroWriteRegisterEnable[9])
						Reg0[ 72: 79] <= in_ZeroWriteData[ 72: 79];
					if (in_ZeroWriteRegisterEnable[10])
						Reg0[ 80: 87] <= in_ZeroWriteData[ 80: 87];
					if (in_ZeroWriteRegisterEnable[11])
						Reg0[ 88: 95] <= in_ZeroWriteData[ 88: 95];
					if (in_ZeroWriteRegisterEnable[12])
						Reg0[ 96:103] <= in_ZeroWriteData[ 96:103];
					if (in_ZeroWriteRegisterEnable[13])
						Reg0[104:111] <= in_ZeroWriteData[104:111];
					if (in_ZeroWriteRegisterEnable[14])
						Reg0[112:119] <= in_ZeroWriteData[112:119];
					if (in_ZeroWriteRegisterEnable[15])
						Reg0[120:127] <= in_ZeroWriteData[120:127];
				  end
      6'b010000 : Reg0 <= in_FirstWriteData;
      6'b001000 : Reg0 <= in_SecondWriteData;
      6'b000100 : Reg0 <= in_ThirdWriteData;
      6'b000010 : Reg0 <= in_FourthWriteData;
      6'b000001 : Reg0 <= in_FifthWriteData;
      default   : Reg0 <= Reg0;
    endcase
  end
  else
  begin
    Reg0 <= Reg0;
  end
end
//write Reg1
always @ ( posedge clk or negedge rst_n )
begin
  if( !rst_n )
  begin
    Reg1 <= 128'h0;
  end
  else if ( | Reg1WriteMask )
  begin
    case ( Reg1WriteMask )
      6'b100000 : begin
					if (in_ZeroWriteRegisterEnable[0])
						Reg1[  0:  7] <= in_ZeroWriteData[  0:  7];
					if (in_ZeroWriteRegisterEnable[1])
						Reg1[  8: 15] <= in_ZeroWriteData[  8: 15];
					if (in_ZeroWriteRegisterEnable[2])
						Reg1[ 16: 23] <= in_ZeroWriteData[ 16: 23];
					if (in_ZeroWriteRegisterEnable[3])
						Reg1[ 24: 31] <= in_ZeroWriteData[ 24: 31];
					if (in_ZeroWriteRegisterEnable[4])
						Reg1[ 32: 39] <= in_ZeroWriteData[ 32: 39];
					if (in_ZeroWriteRegisterEnable[5])
						Reg1[ 40: 47] <= in_ZeroWriteData[ 40: 47];
					if (in_ZeroWriteRegisterEnable[6])
						Reg1[ 48: 55] <= in_ZeroWriteData[ 48: 55];
					if (in_ZeroWriteRegisterEnable[7])
						Reg1[ 56: 63] <= in_ZeroWriteData[ 56: 63];
					if (in_ZeroWriteRegisterEnable[8])
						Reg1[ 64: 71] <= in_ZeroWriteData[ 64: 71];
					if (in_ZeroWriteRegisterEnable[9])
						Reg1[ 72: 79] <= in_ZeroWriteData[ 72: 79];
					if (in_ZeroWriteRegisterEnable[10])
						Reg1[ 80: 87] <= in_ZeroWriteData[ 80: 87];
					if (in_ZeroWriteRegisterEnable[11])
						Reg1[ 88: 95] <= in_ZeroWriteData[ 88: 95];
					if (in_ZeroWriteRegisterEnable[12])
						Reg1[ 96:103] <= in_ZeroWriteData[ 96:103];
					if (in_ZeroWriteRegisterEnable[13])
						Reg1[104:111] <= in_ZeroWriteData[104:111];
					if (in_ZeroWriteRegisterEnable[14])
						Reg1[112:119] <= in_ZeroWriteData[112:119];
					if (in_ZeroWriteRegisterEnable[15])
						Reg1[120:127] <= in_ZeroWriteData[120:127];
				  end
      6'b010000 : Reg1 <= in_FirstWriteData;
      6'b001000 : Reg1 <= in_SecondWriteData;
      6'b000100 : Reg1 <= in_ThirdWriteData;
      6'b000010 : Reg1 <= in_FourthWriteData;
      6'b000001 : Reg1 <= in_FifthWriteData;
      default   : Reg1 <= Reg1;
    endcase
  end
  else
  begin
    Reg1 <= Reg1;
  end
end
//write Reg2
always @ ( posedge clk or negedge rst_n )
begin
  if( !rst_n )
  begin
    Reg2 <= 128'h0;
  end
  else if ( | Reg2WriteMask )
  begin
    case ( Reg2WriteMask )
      6'b100000 : begin
					if (in_ZeroWriteRegisterEnable[0])
						Reg2[  0:  7] <= in_ZeroWriteData[  0:  7];
					if (in_ZeroWriteRegisterEnable[1])
						Reg2[  8: 15] <= in_ZeroWriteData[  8: 15];
					if (in_ZeroWriteRegisterEnable[2])
						Reg2[ 16: 23] <= in_ZeroWriteData[ 16: 23];
					if (in_ZeroWriteRegisterEnable[3])
						Reg2[ 24: 31] <= in_ZeroWriteData[ 24: 31];
					if (in_ZeroWriteRegisterEnable[4])
						Reg2[ 32: 39] <= in_ZeroWriteData[ 32: 39];
					if (in_ZeroWriteRegisterEnable[5])
						Reg2[ 40: 47] <= in_ZeroWriteData[ 40: 47];
					if (in_ZeroWriteRegisterEnable[6])
						Reg2[ 48: 55] <= in_ZeroWriteData[ 48: 55];
					if (in_ZeroWriteRegisterEnable[7])
						Reg2[ 56: 63] <= in_ZeroWriteData[ 56: 63];
					if (in_ZeroWriteRegisterEnable[8])
						Reg2[ 64: 71] <= in_ZeroWriteData[ 64: 71];
					if (in_ZeroWriteRegisterEnable[9])
						Reg2[ 72: 79] <= in_ZeroWriteData[ 72: 79];
					if (in_ZeroWriteRegisterEnable[10])
						Reg2[ 80: 87] <= in_ZeroWriteData[ 80: 87];
					if (in_ZeroWriteRegisterEnable[11])
						Reg2[ 88: 95] <= in_ZeroWriteData[ 88: 95];
					if (in_ZeroWriteRegisterEnable[12])
						Reg2[ 96:103] <= in_ZeroWriteData[ 96:103];
					if (in_ZeroWriteRegisterEnable[13])
						Reg2[104:111] <= in_ZeroWriteData[104:111];
					if (in_ZeroWriteRegisterEnable[14])
						Reg2[112:119] <= in_ZeroWriteData[112:119];
					if (in_ZeroWriteRegisterEnable[15])
						Reg2[120:127] <= in_ZeroWriteData[120:127];
				  end
      6'b010000 : Reg2 <= in_FirstWriteData;
      6'b001000 : Reg2 <= in_SecondWriteData;
      6'b000100 : Reg2 <= in_ThirdWriteData;
      6'b000010 : Reg2 <= in_FourthWriteData;
      6'b000001 : Reg2 <= in_FifthWriteData;
      default   : Reg2 <= Reg2;
    endcase
  end
  else
  begin
    Reg2 <= Reg2;
  end
end
//write Reg3
always @ ( posedge clk or negedge rst_n )
begin
  if( !rst_n )
  begin
    Reg3 <= 128'h0;
  end
  else if ( | Reg3WriteMask )
  begin
    case ( Reg3WriteMask )
      6'b100000 : begin
					if (in_ZeroWriteRegisterEnable[0])
						Reg3[  0:  7] <= in_ZeroWriteData[  0:  7];
					if (in_ZeroWriteRegisterEnable[1])
						Reg3[  8: 15] <= in_ZeroWriteData[  8: 15];
					if (in_ZeroWriteRegisterEnable[2])
						Reg3[ 16: 23] <= in_ZeroWriteData[ 16: 23];
					if (in_ZeroWriteRegisterEnable[3])
						Reg3[ 24: 31] <= in_ZeroWriteData[ 24: 31];
					if (in_ZeroWriteRegisterEnable[4])
						Reg3[ 32: 39] <= in_ZeroWriteData[ 32: 39];
					if (in_ZeroWriteRegisterEnable[5])
						Reg3[ 40: 47] <= in_ZeroWriteData[ 40: 47];
					if (in_ZeroWriteRegisterEnable[6])
						Reg3[ 48: 55] <= in_ZeroWriteData[ 48: 55];
					if (in_ZeroWriteRegisterEnable[7])
						Reg3[ 56: 63] <= in_ZeroWriteData[ 56: 63];
					if (in_ZeroWriteRegisterEnable[8])
						Reg3[ 64: 71] <= in_ZeroWriteData[ 64: 71];
					if (in_ZeroWriteRegisterEnable[9])
						Reg3[ 72: 79] <= in_ZeroWriteData[ 72: 79];
					if (in_ZeroWriteRegisterEnable[10])
						Reg3[ 80: 87] <= in_ZeroWriteData[ 80: 87];
					if (in_ZeroWriteRegisterEnable[11])
						Reg3[ 88: 95] <= in_ZeroWriteData[ 88: 95];
					if (in_ZeroWriteRegisterEnable[12])
						Reg3[ 96:103] <= in_ZeroWriteData[ 96:103];
					if (in_ZeroWriteRegisterEnable[13])
						Reg3[104:111] <= in_ZeroWriteData[104:111];
					if (in_ZeroWriteRegisterEnable[14])
						Reg3[112:119] <= in_ZeroWriteData[112:119];
					if (in_ZeroWriteRegisterEnable[15])
						Reg3[120:127] <= in_ZeroWriteData[120:127];
				  end
      6'b010000 : Reg3 <= in_FirstWriteData;
      6'b001000 : Reg3 <= in_SecondWriteData;
      6'b000100 : Reg3 <= in_ThirdWriteData;
      6'b000010 : Reg3 <= in_FourthWriteData;
      6'b000001 : Reg3 <= in_FifthWriteData;
      default   : Reg3 <= Reg3;
    endcase
  end
  else
  begin
    Reg3 <= Reg3;
  end
end
//write Reg4
always @ ( posedge clk or negedge rst_n )
begin
  if( !rst_n )
  begin
    Reg4 <= 128'h0;
  end
  else if ( | Reg4WriteMask )
  begin
    case ( Reg4WriteMask )
      6'b100000 : begin
					if (in_ZeroWriteRegisterEnable[0])
						Reg4[  0:  7] <= in_ZeroWriteData[  0:  7];
					if (in_ZeroWriteRegisterEnable[1])
						Reg4[  8: 15] <= in_ZeroWriteData[  8: 15];
					if (in_ZeroWriteRegisterEnable[2])
						Reg4[ 16: 23] <= in_ZeroWriteData[ 16: 23];
					if (in_ZeroWriteRegisterEnable[3])
						Reg4[ 24: 31] <= in_ZeroWriteData[ 24: 31];
					if (in_ZeroWriteRegisterEnable[4])
						Reg4[ 32: 39] <= in_ZeroWriteData[ 32: 39];
					if (in_ZeroWriteRegisterEnable[5])
						Reg4[ 40: 47] <= in_ZeroWriteData[ 40: 47];
					if (in_ZeroWriteRegisterEnable[6])
						Reg4[ 48: 55] <= in_ZeroWriteData[ 48: 55];
					if (in_ZeroWriteRegisterEnable[7])
						Reg4[ 56: 63] <= in_ZeroWriteData[ 56: 63];
					if (in_ZeroWriteRegisterEnable[8])
						Reg4[ 64: 71] <= in_ZeroWriteData[ 64: 71];
					if (in_ZeroWriteRegisterEnable[9])
						Reg4[ 72: 79] <= in_ZeroWriteData[ 72: 79];
					if (in_ZeroWriteRegisterEnable[10])
						Reg4[ 80: 87] <= in_ZeroWriteData[ 80: 87];
					if (in_ZeroWriteRegisterEnable[11])
						Reg4[ 88: 95] <= in_ZeroWriteData[ 88: 95];
					if (in_ZeroWriteRegisterEnable[12])
						Reg4[ 96:103] <= in_ZeroWriteData[ 96:103];
					if (in_ZeroWriteRegisterEnable[13])
						Reg4[104:111] <= in_ZeroWriteData[104:111];
					if (in_ZeroWriteRegisterEnable[14])
						Reg4[112:119] <= in_ZeroWriteData[112:119];
					if (in_ZeroWriteRegisterEnable[15])
						Reg4[120:127] <= in_ZeroWriteData[120:127];
				  end
      6'b010000 : Reg4 <= in_FirstWriteData;
      6'b001000 : Reg4 <= in_SecondWriteData;
      6'b000100 : Reg4 <= in_ThirdWriteData;
      6'b000010 : Reg4 <= in_FourthWriteData;
      6'b000001 : Reg4 <= in_FifthWriteData;
      default   : Reg4 <= Reg4;
    endcase
  end
  else
  begin
    Reg4 <= Reg4;
  end
end
//write Reg5
always @ ( posedge clk or negedge rst_n )
begin
  if( !rst_n )
  begin
    Reg5 <= 128'h0;
  end
  else if ( | Reg5WriteMask )
  begin
    case ( Reg5WriteMask )
      6'b100000 : begin
					if (in_ZeroWriteRegisterEnable[0])
						Reg5[  0:  7] <= in_ZeroWriteData[  0:  7];
					if (in_ZeroWriteRegisterEnable[1])
						Reg5[  8: 15] <= in_ZeroWriteData[  8: 15];
					if (in_ZeroWriteRegisterEnable[2])
						Reg5[ 16: 23] <= in_ZeroWriteData[ 16: 23];
					if (in_ZeroWriteRegisterEnable[3])
						Reg5[ 24: 31] <= in_ZeroWriteData[ 24: 31];
					if (in_ZeroWriteRegisterEnable[4])
						Reg5[ 32: 39] <= in_ZeroWriteData[ 32: 39];
					if (in_ZeroWriteRegisterEnable[5])
						Reg5[ 40: 47] <= in_ZeroWriteData[ 40: 47];
					if (in_ZeroWriteRegisterEnable[6])
						Reg5[ 48: 55] <= in_ZeroWriteData[ 48: 55];
					if (in_ZeroWriteRegisterEnable[7])
						Reg5[ 56: 63] <= in_ZeroWriteData[ 56: 63];
					if (in_ZeroWriteRegisterEnable[8])
						Reg5[ 64: 71] <= in_ZeroWriteData[ 64: 71];
					if (in_ZeroWriteRegisterEnable[9])
						Reg5[ 72: 79] <= in_ZeroWriteData[ 72: 79];
					if (in_ZeroWriteRegisterEnable[10])
						Reg5[ 80: 87] <= in_ZeroWriteData[ 80: 87];
					if (in_ZeroWriteRegisterEnable[11])
						Reg5[ 88: 95] <= in_ZeroWriteData[ 88: 95];
					if (in_ZeroWriteRegisterEnable[12])
						Reg5[ 96:103] <= in_ZeroWriteData[ 96:103];
					if (in_ZeroWriteRegisterEnable[13])
						Reg5[104:111] <= in_ZeroWriteData[104:111];
					if (in_ZeroWriteRegisterEnable[14])
						Reg5[112:119] <= in_ZeroWriteData[112:119];
					if (in_ZeroWriteRegisterEnable[15])
						Reg5[120:127] <= in_ZeroWriteData[120:127];
				  end
      6'b010000 : Reg5 <= in_FirstWriteData;
      6'b001000 : Reg5 <= in_SecondWriteData;
      6'b000100 : Reg5 <= in_ThirdWriteData;
      6'b000010 : Reg5 <= in_FourthWriteData;
      6'b000001 : Reg5 <= in_FifthWriteData;
      default   : Reg5 <= Reg5;
    endcase
  end
  else
  begin
    Reg5 <= Reg5;
  end
end
//write Reg6
always @ ( posedge clk or negedge rst_n )
begin
  if( !rst_n )
  begin
    Reg6 <= 128'h0;
  end
  else if ( | Reg6WriteMask )
  begin
    case ( Reg6WriteMask )
      6'b100000 : begin
					if (in_ZeroWriteRegisterEnable[0])
						Reg6[  0:  7] <= in_ZeroWriteData[  0:  7];
					if (in_ZeroWriteRegisterEnable[1])
						Reg6[  8: 15] <= in_ZeroWriteData[  8: 15];
					if (in_ZeroWriteRegisterEnable[2])
						Reg6[ 16: 23] <= in_ZeroWriteData[ 16: 23];
					if (in_ZeroWriteRegisterEnable[3])
						Reg6[ 24: 31] <= in_ZeroWriteData[ 24: 31];
					if (in_ZeroWriteRegisterEnable[4])
						Reg6[ 32: 39] <= in_ZeroWriteData[ 32: 39];
					if (in_ZeroWriteRegisterEnable[5])
						Reg6[ 40: 47] <= in_ZeroWriteData[ 40: 47];
					if (in_ZeroWriteRegisterEnable[6])
						Reg6[ 48: 55] <= in_ZeroWriteData[ 48: 55];
					if (in_ZeroWriteRegisterEnable[7])
						Reg6[ 56: 63] <= in_ZeroWriteData[ 56: 63];
					if (in_ZeroWriteRegisterEnable[8])
						Reg6[ 64: 71] <= in_ZeroWriteData[ 64: 71];
					if (in_ZeroWriteRegisterEnable[9])
						Reg6[ 72: 79] <= in_ZeroWriteData[ 72: 79];
					if (in_ZeroWriteRegisterEnable[10])
						Reg6[ 80: 87] <= in_ZeroWriteData[ 80: 87];
					if (in_ZeroWriteRegisterEnable[11])
						Reg6[ 88: 95] <= in_ZeroWriteData[ 88: 95];
					if (in_ZeroWriteRegisterEnable[12])
						Reg6[ 96:103] <= in_ZeroWriteData[ 96:103];
					if (in_ZeroWriteRegisterEnable[13])
						Reg6[104:111] <= in_ZeroWriteData[104:111];
					if (in_ZeroWriteRegisterEnable[14])
						Reg6[112:119] <= in_ZeroWriteData[112:119];
					if (in_ZeroWriteRegisterEnable[15])
						Reg6[120:127] <= in_ZeroWriteData[120:127];
				  end
      6'b010000 : Reg6 <= in_FirstWriteData;
      6'b001000 : Reg6 <= in_SecondWriteData;
      6'b000100 : Reg6 <= in_ThirdWriteData;
      6'b000010 : Reg6 <= in_FourthWriteData;
      6'b000001 : Reg6 <= in_FifthWriteData;
      default   : Reg6 <= Reg6;
    endcase
  end
  else
  begin
    Reg6 <= Reg6;
  end
end
//write Reg7
always @ ( posedge clk or negedge rst_n )
begin
  if( !rst_n )
  begin
    Reg7 <= 128'h0;
  end
  else if ( | Reg7WriteMask )
  begin
    case ( Reg7WriteMask )
      6'b100000 : begin
					if (in_ZeroWriteRegisterEnable[0])
						Reg7[  0:  7] <= in_ZeroWriteData[  0:  7];
					if (in_ZeroWriteRegisterEnable[1])
						Reg7[  8: 15] <= in_ZeroWriteData[  8: 15];
					if (in_ZeroWriteRegisterEnable[2])
						Reg7[ 16: 23] <= in_ZeroWriteData[ 16: 23];
					if (in_ZeroWriteRegisterEnable[3])
						Reg7[ 24: 31] <= in_ZeroWriteData[ 24: 31];
					if (in_ZeroWriteRegisterEnable[4])
						Reg7[ 32: 39] <= in_ZeroWriteData[ 32: 39];
					if (in_ZeroWriteRegisterEnable[5])
						Reg7[ 40: 47] <= in_ZeroWriteData[ 40: 47];
					if (in_ZeroWriteRegisterEnable[6])
						Reg7[ 48: 55] <= in_ZeroWriteData[ 48: 55];
					if (in_ZeroWriteRegisterEnable[7])
						Reg7[ 56: 63] <= in_ZeroWriteData[ 56: 63];
					if (in_ZeroWriteRegisterEnable[8])
						Reg7[ 64: 71] <= in_ZeroWriteData[ 64: 71];
					if (in_ZeroWriteRegisterEnable[9])
						Reg7[ 72: 79] <= in_ZeroWriteData[ 72: 79];
					if (in_ZeroWriteRegisterEnable[10])
						Reg7[ 80: 87] <= in_ZeroWriteData[ 80: 87];
					if (in_ZeroWriteRegisterEnable[11])
						Reg7[ 88: 95] <= in_ZeroWriteData[ 88: 95];
					if (in_ZeroWriteRegisterEnable[12])
						Reg7[ 96:103] <= in_ZeroWriteData[ 96:103];
					if (in_ZeroWriteRegisterEnable[13])
						Reg7[104:111] <= in_ZeroWriteData[104:111];
					if (in_ZeroWriteRegisterEnable[14])
						Reg7[112:119] <= in_ZeroWriteData[112:119];
					if (in_ZeroWriteRegisterEnable[15])
						Reg7[120:127] <= in_ZeroWriteData[120:127];
				  end
      6'b010000 : Reg7 <= in_FirstWriteData;
      6'b001000 : Reg7 <= in_SecondWriteData;
      6'b000100 : Reg7 <= in_ThirdWriteData;
      6'b000010 : Reg7 <= in_FourthWriteData;
      6'b000001 : Reg7 <= in_FifthWriteData;
      default   : Reg7 <= Reg7;
    endcase
  end
  else
  begin
    Reg7 <= Reg7;
  end
end
//write Reg8
always @ ( posedge clk or negedge rst_n )
begin
  if( !rst_n )
  begin
    Reg8 <= 128'h0;
  end
  else if ( | Reg8WriteMask )
  begin
    case ( Reg8WriteMask )
      6'b100000 : begin
					if (in_ZeroWriteRegisterEnable[0])
						Reg8[  0:  7] <= in_ZeroWriteData[  0:  7];
					if (in_ZeroWriteRegisterEnable[1])
						Reg8[  8: 15] <= in_ZeroWriteData[  8: 15];
					if (in_ZeroWriteRegisterEnable[2])
						Reg8[ 16: 23] <= in_ZeroWriteData[ 16: 23];
					if (in_ZeroWriteRegisterEnable[3])
						Reg8[ 24: 31] <= in_ZeroWriteData[ 24: 31];
					if (in_ZeroWriteRegisterEnable[4])
						Reg8[ 32: 39] <= in_ZeroWriteData[ 32: 39];
					if (in_ZeroWriteRegisterEnable[5])
						Reg8[ 40: 47] <= in_ZeroWriteData[ 40: 47];
					if (in_ZeroWriteRegisterEnable[6])
						Reg8[ 48: 55] <= in_ZeroWriteData[ 48: 55];
					if (in_ZeroWriteRegisterEnable[7])
						Reg8[ 56: 63] <= in_ZeroWriteData[ 56: 63];
					if (in_ZeroWriteRegisterEnable[8])
						Reg8[ 64: 71] <= in_ZeroWriteData[ 64: 71];
					if (in_ZeroWriteRegisterEnable[9])
						Reg8[ 72: 79] <= in_ZeroWriteData[ 72: 79];
					if (in_ZeroWriteRegisterEnable[10])
						Reg8[ 80: 87] <= in_ZeroWriteData[ 80: 87];
					if (in_ZeroWriteRegisterEnable[11])
						Reg8[ 88: 95] <= in_ZeroWriteData[ 88: 95];
					if (in_ZeroWriteRegisterEnable[12])
						Reg8[ 96:103] <= in_ZeroWriteData[ 96:103];
					if (in_ZeroWriteRegisterEnable[13])
						Reg8[104:111] <= in_ZeroWriteData[104:111];
					if (in_ZeroWriteRegisterEnable[14])
						Reg8[112:119] <= in_ZeroWriteData[112:119];
					if (in_ZeroWriteRegisterEnable[15])
						Reg8[120:127] <= in_ZeroWriteData[120:127];
				  end
      6'b010000 : Reg8 <= in_FirstWriteData;
      6'b001000 : Reg8 <= in_SecondWriteData;
      6'b000100 : Reg8 <= in_ThirdWriteData;
      6'b000010 : Reg8 <= in_FourthWriteData;
      6'b000001 : Reg8 <= in_FifthWriteData;
      default   : Reg8 <= Reg8;
    endcase
  end
  else
  begin
    Reg8 <= Reg8;
  end
end
//write Reg9
always @ ( posedge clk or negedge rst_n )
begin
  if( !rst_n )
  begin
    Reg9 <= 128'h0;
  end
  else if ( | Reg9WriteMask )
  begin
    case ( Reg9WriteMask )
      6'b100000 : begin
					if (in_ZeroWriteRegisterEnable[0])
						Reg9[  0:  7] <= in_ZeroWriteData[  0:  7];
					if (in_ZeroWriteRegisterEnable[1])
						Reg9[  8: 15] <= in_ZeroWriteData[  8: 15];
					if (in_ZeroWriteRegisterEnable[2])
						Reg9[ 16: 23] <= in_ZeroWriteData[ 16: 23];
					if (in_ZeroWriteRegisterEnable[3])
						Reg9[ 24: 31] <= in_ZeroWriteData[ 24: 31];
					if (in_ZeroWriteRegisterEnable[4])
						Reg9[ 32: 39] <= in_ZeroWriteData[ 32: 39];
					if (in_ZeroWriteRegisterEnable[5])
						Reg9[ 40: 47] <= in_ZeroWriteData[ 40: 47];
					if (in_ZeroWriteRegisterEnable[6])
						Reg9[ 48: 55] <= in_ZeroWriteData[ 48: 55];
					if (in_ZeroWriteRegisterEnable[7])
						Reg9[ 56: 63] <= in_ZeroWriteData[ 56: 63];
					if (in_ZeroWriteRegisterEnable[8])
						Reg9[ 64: 71] <= in_ZeroWriteData[ 64: 71];
					if (in_ZeroWriteRegisterEnable[9])
						Reg9[ 72: 79] <= in_ZeroWriteData[ 72: 79];
					if (in_ZeroWriteRegisterEnable[10])
						Reg9[ 80: 87] <= in_ZeroWriteData[ 80: 87];
					if (in_ZeroWriteRegisterEnable[11])
						Reg9[ 88: 95] <= in_ZeroWriteData[ 88: 95];
					if (in_ZeroWriteRegisterEnable[12])
						Reg9[ 96:103] <= in_ZeroWriteData[ 96:103];
					if (in_ZeroWriteRegisterEnable[13])
						Reg9[104:111] <= in_ZeroWriteData[104:111];
					if (in_ZeroWriteRegisterEnable[14])
						Reg9[112:119] <= in_ZeroWriteData[112:119];
					if (in_ZeroWriteRegisterEnable[15])
						Reg9[120:127] <= in_ZeroWriteData[120:127];
				  end
      6'b010000 : Reg9 <= in_FirstWriteData;
      6'b001000 : Reg9 <= in_SecondWriteData;
      6'b000100 : Reg9 <= in_ThirdWriteData;
      6'b000010 : Reg9 <= in_FourthWriteData;
      6'b000001 : Reg9 <= in_FifthWriteData;
      default   : Reg9 <= Reg9;
    endcase
  end
  else
  begin
    Reg9 <= Reg9;
  end
end
//write Reg10
always @ ( posedge clk or negedge rst_n )
begin
  if( !rst_n )
  begin
    Reg10 <= 128'h0;
  end
  else if ( | Reg10WriteMask )
  begin
    case ( Reg10WriteMask )
      6'b100000 : begin
					if (in_ZeroWriteRegisterEnable[0])
						Reg10[  0:  7] <= in_ZeroWriteData[  0:  7];
					if (in_ZeroWriteRegisterEnable[1])
						Reg10[  8: 15] <= in_ZeroWriteData[  8: 15];
					if (in_ZeroWriteRegisterEnable[2])
						Reg10[ 16: 23] <= in_ZeroWriteData[ 16: 23];
					if (in_ZeroWriteRegisterEnable[3])
						Reg10[ 24: 31] <= in_ZeroWriteData[ 24: 31];
					if (in_ZeroWriteRegisterEnable[4])
						Reg10[ 32: 39] <= in_ZeroWriteData[ 32: 39];
					if (in_ZeroWriteRegisterEnable[5])
						Reg10[ 40: 47] <= in_ZeroWriteData[ 40: 47];
					if (in_ZeroWriteRegisterEnable[6])
						Reg10[ 48: 55] <= in_ZeroWriteData[ 48: 55];
					if (in_ZeroWriteRegisterEnable[7])
						Reg10[ 56: 63] <= in_ZeroWriteData[ 56: 63];
					if (in_ZeroWriteRegisterEnable[8])
						Reg10[ 64: 71] <= in_ZeroWriteData[ 64: 71];
					if (in_ZeroWriteRegisterEnable[9])
						Reg10[ 72: 79] <= in_ZeroWriteData[ 72: 79];
					if (in_ZeroWriteRegisterEnable[10])
						Reg10[ 80: 87] <= in_ZeroWriteData[ 80: 87];
					if (in_ZeroWriteRegisterEnable[11])
						Reg10[ 88: 95] <= in_ZeroWriteData[ 88: 95];
					if (in_ZeroWriteRegisterEnable[12])
						Reg10[ 96:103] <= in_ZeroWriteData[ 96:103];
					if (in_ZeroWriteRegisterEnable[13])
						Reg10[104:111] <= in_ZeroWriteData[104:111];
					if (in_ZeroWriteRegisterEnable[14])
						Reg10[112:119] <= in_ZeroWriteData[112:119];
					if (in_ZeroWriteRegisterEnable[15])
						Reg10[120:127] <= in_ZeroWriteData[120:127];
				  end
      6'b010000 : Reg10 <= in_FirstWriteData;
      6'b001000 : Reg10 <= in_SecondWriteData;
      6'b000100 : Reg10 <= in_ThirdWriteData;
      6'b000010 : Reg10 <= in_FourthWriteData;
      6'b000001 : Reg10 <= in_FifthWriteData;
      default   : Reg10 <= Reg10;
    endcase
  end
  else
  begin
    Reg10 <= Reg10;
  end
end
//write Reg11
always @ ( posedge clk or negedge rst_n )
begin
  if( !rst_n )
  begin
    Reg11 <= 128'h0;
  end
  else if ( | Reg11WriteMask )
  begin
    case ( Reg11WriteMask )
      6'b100000 : begin
					if (in_ZeroWriteRegisterEnable[0])
						Reg11[  0:  7] <= in_ZeroWriteData[  0:  7];
					if (in_ZeroWriteRegisterEnable[1])
						Reg11[  8: 15] <= in_ZeroWriteData[  8: 15];
					if (in_ZeroWriteRegisterEnable[2])
						Reg11[ 16: 23] <= in_ZeroWriteData[ 16: 23];
					if (in_ZeroWriteRegisterEnable[3])
						Reg11[ 24: 31] <= in_ZeroWriteData[ 24: 31];
					if (in_ZeroWriteRegisterEnable[4])
						Reg11[ 32: 39] <= in_ZeroWriteData[ 32: 39];
					if (in_ZeroWriteRegisterEnable[5])
						Reg11[ 40: 47] <= in_ZeroWriteData[ 40: 47];
					if (in_ZeroWriteRegisterEnable[6])
						Reg11[ 48: 55] <= in_ZeroWriteData[ 48: 55];
					if (in_ZeroWriteRegisterEnable[7])
						Reg11[ 56: 63] <= in_ZeroWriteData[ 56: 63];
					if (in_ZeroWriteRegisterEnable[8])
						Reg11[ 64: 71] <= in_ZeroWriteData[ 64: 71];
					if (in_ZeroWriteRegisterEnable[9])
						Reg11[ 72: 79] <= in_ZeroWriteData[ 72: 79];
					if (in_ZeroWriteRegisterEnable[10])
						Reg11[ 80: 87] <= in_ZeroWriteData[ 80: 87];
					if (in_ZeroWriteRegisterEnable[11])
						Reg11[ 88: 95] <= in_ZeroWriteData[ 88: 95];
					if (in_ZeroWriteRegisterEnable[12])
						Reg11[ 96:103] <= in_ZeroWriteData[ 96:103];
					if (in_ZeroWriteRegisterEnable[13])
						Reg11[104:111] <= in_ZeroWriteData[104:111];
					if (in_ZeroWriteRegisterEnable[14])
						Reg11[112:119] <= in_ZeroWriteData[112:119];
					if (in_ZeroWriteRegisterEnable[15])
						Reg11[120:127] <= in_ZeroWriteData[120:127];
				  end
      6'b010000 : Reg11 <= in_FirstWriteData;
      6'b001000 : Reg11 <= in_SecondWriteData;
      6'b000100 : Reg11 <= in_ThirdWriteData;
      6'b000010 : Reg11 <= in_FourthWriteData;
      6'b000001 : Reg11 <= in_FifthWriteData;
      default   : Reg11 <= Reg11;
    endcase
  end
  else
  begin
    Reg11 <= Reg11;
  end
end
//write Reg12
always @ ( posedge clk or negedge rst_n )
begin
  if( !rst_n )
  begin
    Reg12 <= 128'h0;
  end
  else if ( | Reg12WriteMask )
  begin
    case ( Reg12WriteMask )
      6'b100000 : begin
					if (in_ZeroWriteRegisterEnable[0])
						Reg12[  0:  7] <= in_ZeroWriteData[  0:  7];
					if (in_ZeroWriteRegisterEnable[1])
						Reg12[  8: 15] <= in_ZeroWriteData[  8: 15];
					if (in_ZeroWriteRegisterEnable[2])
						Reg12[ 16: 23] <= in_ZeroWriteData[ 16: 23];
					if (in_ZeroWriteRegisterEnable[3])
						Reg12[ 24: 31] <= in_ZeroWriteData[ 24: 31];
					if (in_ZeroWriteRegisterEnable[4])
						Reg12[ 32: 39] <= in_ZeroWriteData[ 32: 39];
					if (in_ZeroWriteRegisterEnable[5])
						Reg12[ 40: 47] <= in_ZeroWriteData[ 40: 47];
					if (in_ZeroWriteRegisterEnable[6])
						Reg12[ 48: 55] <= in_ZeroWriteData[ 48: 55];
					if (in_ZeroWriteRegisterEnable[7])
						Reg12[ 56: 63] <= in_ZeroWriteData[ 56: 63];
					if (in_ZeroWriteRegisterEnable[8])
						Reg12[ 64: 71] <= in_ZeroWriteData[ 64: 71];
					if (in_ZeroWriteRegisterEnable[9])
						Reg12[ 72: 79] <= in_ZeroWriteData[ 72: 79];
					if (in_ZeroWriteRegisterEnable[10])
						Reg12[ 80: 87] <= in_ZeroWriteData[ 80: 87];
					if (in_ZeroWriteRegisterEnable[11])
						Reg12[ 88: 95] <= in_ZeroWriteData[ 88: 95];
					if (in_ZeroWriteRegisterEnable[12])
						Reg12[ 96:103] <= in_ZeroWriteData[ 96:103];
					if (in_ZeroWriteRegisterEnable[13])
						Reg12[104:111] <= in_ZeroWriteData[104:111];
					if (in_ZeroWriteRegisterEnable[14])
						Reg12[112:119] <= in_ZeroWriteData[112:119];
					if (in_ZeroWriteRegisterEnable[15])
						Reg12[120:127] <= in_ZeroWriteData[120:127];
				  end
      6'b010000 : Reg12 <= in_FirstWriteData;
      6'b001000 : Reg12 <= in_SecondWriteData;
      6'b000100 : Reg12 <= in_ThirdWriteData;
      6'b000010 : Reg12 <= in_FourthWriteData;
      6'b000001 : Reg12 <= in_FifthWriteData;
      default   : Reg12 <= Reg12;
    endcase
  end
  else
  begin
    Reg12 <= Reg12;
  end
end
//write Reg13
always @ ( posedge clk or negedge rst_n )
begin
  if( !rst_n )
  begin
    Reg13 <= 128'h0;
  end
  else if ( | Reg13WriteMask )
  begin
    case ( Reg13WriteMask )
      6'b100000 : begin
					if (in_ZeroWriteRegisterEnable[0])
						Reg13[  0:  7] <= in_ZeroWriteData[  0:  7];
					if (in_ZeroWriteRegisterEnable[1])
						Reg13[  8: 15] <= in_ZeroWriteData[  8: 15];
					if (in_ZeroWriteRegisterEnable[2])
						Reg13[ 16: 23] <= in_ZeroWriteData[ 16: 23];
					if (in_ZeroWriteRegisterEnable[3])
						Reg13[ 24: 31] <= in_ZeroWriteData[ 24: 31];
					if (in_ZeroWriteRegisterEnable[4])
						Reg13[ 32: 39] <= in_ZeroWriteData[ 32: 39];
					if (in_ZeroWriteRegisterEnable[5])
						Reg13[ 40: 47] <= in_ZeroWriteData[ 40: 47];
					if (in_ZeroWriteRegisterEnable[6])
						Reg13[ 48: 55] <= in_ZeroWriteData[ 48: 55];
					if (in_ZeroWriteRegisterEnable[7])
						Reg13[ 56: 63] <= in_ZeroWriteData[ 56: 63];
					if (in_ZeroWriteRegisterEnable[8])
						Reg13[ 64: 71] <= in_ZeroWriteData[ 64: 71];
					if (in_ZeroWriteRegisterEnable[9])
						Reg13[ 72: 79] <= in_ZeroWriteData[ 72: 79];
					if (in_ZeroWriteRegisterEnable[10])
						Reg13[ 80: 87] <= in_ZeroWriteData[ 80: 87];
					if (in_ZeroWriteRegisterEnable[11])
						Reg13[ 88: 95] <= in_ZeroWriteData[ 88: 95];
					if (in_ZeroWriteRegisterEnable[12])
						Reg13[ 96:103] <= in_ZeroWriteData[ 96:103];
					if (in_ZeroWriteRegisterEnable[13])
						Reg13[104:111] <= in_ZeroWriteData[104:111];
					if (in_ZeroWriteRegisterEnable[14])
						Reg13[112:119] <= in_ZeroWriteData[112:119];
					if (in_ZeroWriteRegisterEnable[15])
						Reg13[120:127] <= in_ZeroWriteData[120:127];
				  end
      6'b010000 : Reg13 <= in_FirstWriteData;
      6'b001000 : Reg13 <= in_SecondWriteData;
      6'b000100 : Reg13 <= in_ThirdWriteData;
      6'b000010 : Reg13 <= in_FourthWriteData;
      6'b000001 : Reg13 <= in_FifthWriteData;
      default   : Reg13 <= Reg13;
    endcase
  end
  else
  begin
    Reg13 <= Reg13;
  end
end
//write Reg14
always @ ( posedge clk or negedge rst_n )
begin
  if( !rst_n )
  begin
    Reg14 <= 128'h0;
  end
  else if ( | Reg14WriteMask )
  begin
    case ( Reg14WriteMask )
      6'b100000 : begin
					if (in_ZeroWriteRegisterEnable[0])
						Reg14[  0:  7] <= in_ZeroWriteData[  0:  7];
					if (in_ZeroWriteRegisterEnable[1])
						Reg14[  8: 15] <= in_ZeroWriteData[  8: 15];
					if (in_ZeroWriteRegisterEnable[2])
						Reg14[ 16: 23] <= in_ZeroWriteData[ 16: 23];
					if (in_ZeroWriteRegisterEnable[3])
						Reg14[ 24: 31] <= in_ZeroWriteData[ 24: 31];
					if (in_ZeroWriteRegisterEnable[4])
						Reg14[ 32: 39] <= in_ZeroWriteData[ 32: 39];
					if (in_ZeroWriteRegisterEnable[5])
						Reg14[ 40: 47] <= in_ZeroWriteData[ 40: 47];
					if (in_ZeroWriteRegisterEnable[6])
						Reg14[ 48: 55] <= in_ZeroWriteData[ 48: 55];
					if (in_ZeroWriteRegisterEnable[7])
						Reg14[ 56: 63] <= in_ZeroWriteData[ 56: 63];
					if (in_ZeroWriteRegisterEnable[8])
						Reg14[ 64: 71] <= in_ZeroWriteData[ 64: 71];
					if (in_ZeroWriteRegisterEnable[9])
						Reg14[ 72: 79] <= in_ZeroWriteData[ 72: 79];
					if (in_ZeroWriteRegisterEnable[10])
						Reg14[ 80: 87] <= in_ZeroWriteData[ 80: 87];
					if (in_ZeroWriteRegisterEnable[11])
						Reg14[ 88: 95] <= in_ZeroWriteData[ 88: 95];
					if (in_ZeroWriteRegisterEnable[12])
						Reg14[ 96:103] <= in_ZeroWriteData[ 96:103];
					if (in_ZeroWriteRegisterEnable[13])
						Reg14[104:111] <= in_ZeroWriteData[104:111];
					if (in_ZeroWriteRegisterEnable[14])
						Reg14[112:119] <= in_ZeroWriteData[112:119];
					if (in_ZeroWriteRegisterEnable[15])
						Reg14[120:127] <= in_ZeroWriteData[120:127];
				  end
      6'b010000 : Reg14 <= in_FirstWriteData;
      6'b001000 : Reg14 <= in_SecondWriteData;
      6'b000100 : Reg14 <= in_ThirdWriteData;
      6'b000010 : Reg14 <= in_FourthWriteData;
      6'b000001 : Reg14 <= in_FifthWriteData;
      default   : Reg14 <= Reg14;
    endcase
  end
  else
  begin
    Reg14 <= Reg14;
  end
end
//write Reg15
always @ ( posedge clk or negedge rst_n )
begin
  if( !rst_n )
  begin
    Reg15 <= 128'h0;
  end
  else if ( | Reg15WriteMask )
  begin
    case ( Reg15WriteMask )
      6'b100000 : begin
					if (in_ZeroWriteRegisterEnable[0])
						Reg15[  0:  7] <= in_ZeroWriteData[  0:  7];
					if (in_ZeroWriteRegisterEnable[1])
						Reg15[  8: 15] <= in_ZeroWriteData[  8: 15];
					if (in_ZeroWriteRegisterEnable[2])
						Reg15[ 16: 23] <= in_ZeroWriteData[ 16: 23];
					if (in_ZeroWriteRegisterEnable[3])
						Reg15[ 24: 31] <= in_ZeroWriteData[ 24: 31];
					if (in_ZeroWriteRegisterEnable[4])
						Reg15[ 32: 39] <= in_ZeroWriteData[ 32: 39];
					if (in_ZeroWriteRegisterEnable[5])
						Reg15[ 40: 47] <= in_ZeroWriteData[ 40: 47];
					if (in_ZeroWriteRegisterEnable[6])
						Reg15[ 48: 55] <= in_ZeroWriteData[ 48: 55];
					if (in_ZeroWriteRegisterEnable[7])
						Reg15[ 56: 63] <= in_ZeroWriteData[ 56: 63];
					if (in_ZeroWriteRegisterEnable[8])
						Reg15[ 64: 71] <= in_ZeroWriteData[ 64: 71];
					if (in_ZeroWriteRegisterEnable[9])
						Reg15[ 72: 79] <= in_ZeroWriteData[ 72: 79];
					if (in_ZeroWriteRegisterEnable[10])
						Reg15[ 80: 87] <= in_ZeroWriteData[ 80: 87];
					if (in_ZeroWriteRegisterEnable[11])
						Reg15[ 88: 95] <= in_ZeroWriteData[ 88: 95];
					if (in_ZeroWriteRegisterEnable[12])
						Reg15[ 96:103] <= in_ZeroWriteData[ 96:103];
					if (in_ZeroWriteRegisterEnable[13])
						Reg15[104:111] <= in_ZeroWriteData[104:111];
					if (in_ZeroWriteRegisterEnable[14])
						Reg15[112:119] <= in_ZeroWriteData[112:119];
					if (in_ZeroWriteRegisterEnable[15])
						Reg15[120:127] <= in_ZeroWriteData[120:127];
				  end
      6'b010000 : Reg15 <= in_FirstWriteData;
      6'b001000 : Reg15 <= in_SecondWriteData;
      6'b000100 : Reg15 <= in_ThirdWriteData;
      6'b000010 : Reg15 <= in_FourthWriteData;
      6'b000001 : Reg15 <= in_FifthWriteData;
      default   : Reg15 <= Reg15;
    endcase
  end
  else
  begin
    Reg15 <= Reg15;
  end
end
//write Reg16
always @ ( posedge clk or negedge rst_n )
begin
  if( !rst_n )
  begin
    Reg16 <= 128'h0;
  end
  else if ( | Reg16WriteMask )
  begin
    case ( Reg16WriteMask )
      6'b100000 : begin
					if (in_ZeroWriteRegisterEnable[0])
						Reg16[  0:  7] <= in_ZeroWriteData[  0:  7];
					if (in_ZeroWriteRegisterEnable[1])
						Reg16[  8: 15] <= in_ZeroWriteData[  8: 15];
					if (in_ZeroWriteRegisterEnable[2])
						Reg16[ 16: 23] <= in_ZeroWriteData[ 16: 23];
					if (in_ZeroWriteRegisterEnable[3])
						Reg16[ 24: 31] <= in_ZeroWriteData[ 24: 31];
					if (in_ZeroWriteRegisterEnable[4])
						Reg16[ 32: 39] <= in_ZeroWriteData[ 32: 39];
					if (in_ZeroWriteRegisterEnable[5])
						Reg16[ 40: 47] <= in_ZeroWriteData[ 40: 47];
					if (in_ZeroWriteRegisterEnable[6])
						Reg16[ 48: 55] <= in_ZeroWriteData[ 48: 55];
					if (in_ZeroWriteRegisterEnable[7])
						Reg16[ 56: 63] <= in_ZeroWriteData[ 56: 63];
					if (in_ZeroWriteRegisterEnable[8])
						Reg16[ 64: 71] <= in_ZeroWriteData[ 64: 71];
					if (in_ZeroWriteRegisterEnable[9])
						Reg16[ 72: 79] <= in_ZeroWriteData[ 72: 79];
					if (in_ZeroWriteRegisterEnable[10])
						Reg16[ 80: 87] <= in_ZeroWriteData[ 80: 87];
					if (in_ZeroWriteRegisterEnable[11])
						Reg16[ 88: 95] <= in_ZeroWriteData[ 88: 95];
					if (in_ZeroWriteRegisterEnable[12])
						Reg16[ 96:103] <= in_ZeroWriteData[ 96:103];
					if (in_ZeroWriteRegisterEnable[13])
						Reg16[104:111] <= in_ZeroWriteData[104:111];
					if (in_ZeroWriteRegisterEnable[14])
						Reg16[112:119] <= in_ZeroWriteData[112:119];
					if (in_ZeroWriteRegisterEnable[15])
						Reg16[120:127] <= in_ZeroWriteData[120:127];
				  end
      6'b010000 : Reg16 <= in_FirstWriteData;
      6'b001000 : Reg16 <= in_SecondWriteData;
      6'b000100 : Reg16 <= in_ThirdWriteData;
      6'b000010 : Reg16 <= in_FourthWriteData;
      6'b000001 : Reg16 <= in_FifthWriteData;
      default   : Reg16 <= Reg16;
    endcase
  end
  else
  begin
    Reg16 <= Reg16;
  end
end
//write Reg17
always @ ( posedge clk or negedge rst_n )
begin
  if( !rst_n )
  begin
    Reg17 <= 128'h0;
  end
  else if ( | Reg17WriteMask )
  begin
    case ( Reg17WriteMask )
      6'b100000 : begin
					if (in_ZeroWriteRegisterEnable[0])
						Reg17[  0:  7] <= in_ZeroWriteData[  0:  7];
					if (in_ZeroWriteRegisterEnable[1])
						Reg17[  8: 15] <= in_ZeroWriteData[  8: 15];
					if (in_ZeroWriteRegisterEnable[2])
						Reg17[ 16: 23] <= in_ZeroWriteData[ 16: 23];
					if (in_ZeroWriteRegisterEnable[3])
						Reg17[ 24: 31] <= in_ZeroWriteData[ 24: 31];
					if (in_ZeroWriteRegisterEnable[4])
						Reg17[ 32: 39] <= in_ZeroWriteData[ 32: 39];
					if (in_ZeroWriteRegisterEnable[5])
						Reg17[ 40: 47] <= in_ZeroWriteData[ 40: 47];
					if (in_ZeroWriteRegisterEnable[6])
						Reg17[ 48: 55] <= in_ZeroWriteData[ 48: 55];
					if (in_ZeroWriteRegisterEnable[7])
						Reg17[ 56: 63] <= in_ZeroWriteData[ 56: 63];
					if (in_ZeroWriteRegisterEnable[8])
						Reg17[ 64: 71] <= in_ZeroWriteData[ 64: 71];
					if (in_ZeroWriteRegisterEnable[9])
						Reg17[ 72: 79] <= in_ZeroWriteData[ 72: 79];
					if (in_ZeroWriteRegisterEnable[10])
						Reg17[ 80: 87] <= in_ZeroWriteData[ 80: 87];
					if (in_ZeroWriteRegisterEnable[11])
						Reg17[ 88: 95] <= in_ZeroWriteData[ 88: 95];
					if (in_ZeroWriteRegisterEnable[12])
						Reg17[ 96:103] <= in_ZeroWriteData[ 96:103];
					if (in_ZeroWriteRegisterEnable[13])
						Reg17[104:111] <= in_ZeroWriteData[104:111];
					if (in_ZeroWriteRegisterEnable[14])
						Reg17[112:119] <= in_ZeroWriteData[112:119];
					if (in_ZeroWriteRegisterEnable[15])
						Reg17[120:127] <= in_ZeroWriteData[120:127];
				  end
      6'b010000 : Reg17 <= in_FirstWriteData;
      6'b001000 : Reg17 <= in_SecondWriteData;
      6'b000100 : Reg17 <= in_ThirdWriteData;
      6'b000010 : Reg17 <= in_FourthWriteData;
      6'b000001 : Reg17 <= in_FifthWriteData;
      default   : Reg17 <= Reg17;
    endcase
  end
  else
  begin
    Reg17 <= Reg17;
  end
end
//write Reg18
always @ ( posedge clk or negedge rst_n )
begin
  if( !rst_n )
  begin
    Reg18 <= 128'h0;
  end
  else if ( | Reg18WriteMask )
  begin
    case ( Reg18WriteMask )
      6'b100000 : begin
					if (in_ZeroWriteRegisterEnable[0])
						Reg18[  0:  7] <= in_ZeroWriteData[  0:  7];
					if (in_ZeroWriteRegisterEnable[1])
						Reg18[  8: 15] <= in_ZeroWriteData[  8: 15];
					if (in_ZeroWriteRegisterEnable[2])
						Reg18[ 16: 23] <= in_ZeroWriteData[ 16: 23];
					if (in_ZeroWriteRegisterEnable[3])
						Reg18[ 24: 31] <= in_ZeroWriteData[ 24: 31];
					if (in_ZeroWriteRegisterEnable[4])
						Reg18[ 32: 39] <= in_ZeroWriteData[ 32: 39];
					if (in_ZeroWriteRegisterEnable[5])
						Reg18[ 40: 47] <= in_ZeroWriteData[ 40: 47];
					if (in_ZeroWriteRegisterEnable[6])
						Reg18[ 48: 55] <= in_ZeroWriteData[ 48: 55];
					if (in_ZeroWriteRegisterEnable[7])
						Reg18[ 56: 63] <= in_ZeroWriteData[ 56: 63];
					if (in_ZeroWriteRegisterEnable[8])
						Reg18[ 64: 71] <= in_ZeroWriteData[ 64: 71];
					if (in_ZeroWriteRegisterEnable[9])
						Reg18[ 72: 79] <= in_ZeroWriteData[ 72: 79];
					if (in_ZeroWriteRegisterEnable[10])
						Reg18[ 80: 87] <= in_ZeroWriteData[ 80: 87];
					if (in_ZeroWriteRegisterEnable[11])
						Reg18[ 88: 95] <= in_ZeroWriteData[ 88: 95];
					if (in_ZeroWriteRegisterEnable[12])
						Reg18[ 96:103] <= in_ZeroWriteData[ 96:103];
					if (in_ZeroWriteRegisterEnable[13])
						Reg18[104:111] <= in_ZeroWriteData[104:111];
					if (in_ZeroWriteRegisterEnable[14])
						Reg18[112:119] <= in_ZeroWriteData[112:119];
					if (in_ZeroWriteRegisterEnable[15])
						Reg18[120:127] <= in_ZeroWriteData[120:127];
				  end
      6'b010000 : Reg18 <= in_FirstWriteData;
      6'b001000 : Reg18 <= in_SecondWriteData;
      6'b000100 : Reg18 <= in_ThirdWriteData;
      6'b000010 : Reg18 <= in_FourthWriteData;
      6'b000001 : Reg18 <= in_FifthWriteData;
      default   : Reg18 <= Reg18;
    endcase
  end
  else
  begin
    Reg18 <= Reg18;
  end
end
//write Reg19
always @ ( posedge clk or negedge rst_n )
begin
  if( !rst_n )
  begin
    Reg19 <= 128'h0;
  end
  else if ( | Reg19WriteMask )
  begin
    case ( Reg19WriteMask )
      6'b100000 : begin
					if (in_ZeroWriteRegisterEnable[0])
						Reg19[  0:  7] <= in_ZeroWriteData[  0:  7];
					if (in_ZeroWriteRegisterEnable[1])
						Reg19[  8: 15] <= in_ZeroWriteData[  8: 15];
					if (in_ZeroWriteRegisterEnable[2])
						Reg19[ 16: 23] <= in_ZeroWriteData[ 16: 23];
					if (in_ZeroWriteRegisterEnable[3])
						Reg19[ 24: 31] <= in_ZeroWriteData[ 24: 31];
					if (in_ZeroWriteRegisterEnable[4])
						Reg19[ 32: 39] <= in_ZeroWriteData[ 32: 39];
					if (in_ZeroWriteRegisterEnable[5])
						Reg19[ 40: 47] <= in_ZeroWriteData[ 40: 47];
					if (in_ZeroWriteRegisterEnable[6])
						Reg19[ 48: 55] <= in_ZeroWriteData[ 48: 55];
					if (in_ZeroWriteRegisterEnable[7])
						Reg19[ 56: 63] <= in_ZeroWriteData[ 56: 63];
					if (in_ZeroWriteRegisterEnable[8])
						Reg19[ 64: 71] <= in_ZeroWriteData[ 64: 71];
					if (in_ZeroWriteRegisterEnable[9])
						Reg19[ 72: 79] <= in_ZeroWriteData[ 72: 79];
					if (in_ZeroWriteRegisterEnable[10])
						Reg19[ 80: 87] <= in_ZeroWriteData[ 80: 87];
					if (in_ZeroWriteRegisterEnable[11])
						Reg19[ 88: 95] <= in_ZeroWriteData[ 88: 95];
					if (in_ZeroWriteRegisterEnable[12])
						Reg19[ 96:103] <= in_ZeroWriteData[ 96:103];
					if (in_ZeroWriteRegisterEnable[13])
						Reg19[104:111] <= in_ZeroWriteData[104:111];
					if (in_ZeroWriteRegisterEnable[14])
						Reg19[112:119] <= in_ZeroWriteData[112:119];
					if (in_ZeroWriteRegisterEnable[15])
						Reg19[120:127] <= in_ZeroWriteData[120:127];
				  end
      6'b010000 : Reg19 <= in_FirstWriteData;
      6'b001000 : Reg19 <= in_SecondWriteData;
      6'b000100 : Reg19 <= in_ThirdWriteData;
      6'b000010 : Reg19 <= in_FourthWriteData;
      6'b000001 : Reg19 <= in_FifthWriteData;
      default   : Reg19 <= Reg19;
    endcase
  end
  else
  begin
    Reg19 <= Reg19;
  end
end
//write Reg20
always @ ( posedge clk or negedge rst_n )
begin
  if( !rst_n )
  begin
    Reg20 <= 128'h0;
  end
  else if ( | Reg20WriteMask )
  begin
    case ( Reg20WriteMask )
      6'b100000 : begin
					if (in_ZeroWriteRegisterEnable[0])
						Reg20[  0:  7] <= in_ZeroWriteData[  0:  7];
					if (in_ZeroWriteRegisterEnable[1])
						Reg20[  8: 15] <= in_ZeroWriteData[  8: 15];
					if (in_ZeroWriteRegisterEnable[2])
						Reg20[ 16: 23] <= in_ZeroWriteData[ 16: 23];
					if (in_ZeroWriteRegisterEnable[3])
						Reg20[ 24: 31] <= in_ZeroWriteData[ 24: 31];
					if (in_ZeroWriteRegisterEnable[4])
						Reg20[ 32: 39] <= in_ZeroWriteData[ 32: 39];
					if (in_ZeroWriteRegisterEnable[5])
						Reg20[ 40: 47] <= in_ZeroWriteData[ 40: 47];
					if (in_ZeroWriteRegisterEnable[6])
						Reg20[ 48: 55] <= in_ZeroWriteData[ 48: 55];
					if (in_ZeroWriteRegisterEnable[7])
						Reg20[ 56: 63] <= in_ZeroWriteData[ 56: 63];
					if (in_ZeroWriteRegisterEnable[8])
						Reg20[ 64: 71] <= in_ZeroWriteData[ 64: 71];
					if (in_ZeroWriteRegisterEnable[9])
						Reg20[ 72: 79] <= in_ZeroWriteData[ 72: 79];
					if (in_ZeroWriteRegisterEnable[10])
						Reg20[ 80: 87] <= in_ZeroWriteData[ 80: 87];
					if (in_ZeroWriteRegisterEnable[11])
						Reg20[ 88: 95] <= in_ZeroWriteData[ 88: 95];
					if (in_ZeroWriteRegisterEnable[12])
						Reg20[ 96:103] <= in_ZeroWriteData[ 96:103];
					if (in_ZeroWriteRegisterEnable[13])
						Reg20[104:111] <= in_ZeroWriteData[104:111];
					if (in_ZeroWriteRegisterEnable[14])
						Reg20[112:119] <= in_ZeroWriteData[112:119];
					if (in_ZeroWriteRegisterEnable[15])
						Reg20[120:127] <= in_ZeroWriteData[120:127];
				  end
      6'b010000 : Reg20 <= in_FirstWriteData;
      6'b001000 : Reg20 <= in_SecondWriteData;
      6'b000100 : Reg20 <= in_ThirdWriteData;
      6'b000010 : Reg20 <= in_FourthWriteData;
      6'b000001 : Reg20 <= in_FifthWriteData;
      default   : Reg20 <= Reg20;
    endcase
  end
  else
  begin
    Reg20 <= Reg20;
  end
end
//write Reg21
always @ ( posedge clk or negedge rst_n )
begin
  if( !rst_n )
  begin
    Reg21 <= 128'h0;
  end
  else if ( | Reg21WriteMask )
  begin
    case ( Reg21WriteMask )
      6'b100000 : begin
					if (in_ZeroWriteRegisterEnable[0])
						Reg21[  0:  7] <= in_ZeroWriteData[  0:  7];
					if (in_ZeroWriteRegisterEnable[1])
						Reg21[  8: 15] <= in_ZeroWriteData[  8: 15];
					if (in_ZeroWriteRegisterEnable[2])
						Reg21[ 16: 23] <= in_ZeroWriteData[ 16: 23];
					if (in_ZeroWriteRegisterEnable[3])
						Reg21[ 24: 31] <= in_ZeroWriteData[ 24: 31];
					if (in_ZeroWriteRegisterEnable[4])
						Reg21[ 32: 39] <= in_ZeroWriteData[ 32: 39];
					if (in_ZeroWriteRegisterEnable[5])
						Reg21[ 40: 47] <= in_ZeroWriteData[ 40: 47];
					if (in_ZeroWriteRegisterEnable[6])
						Reg21[ 48: 55] <= in_ZeroWriteData[ 48: 55];
					if (in_ZeroWriteRegisterEnable[7])
						Reg21[ 56: 63] <= in_ZeroWriteData[ 56: 63];
					if (in_ZeroWriteRegisterEnable[8])
						Reg21[ 64: 71] <= in_ZeroWriteData[ 64: 71];
					if (in_ZeroWriteRegisterEnable[9])
						Reg21[ 72: 79] <= in_ZeroWriteData[ 72: 79];
					if (in_ZeroWriteRegisterEnable[10])
						Reg21[ 80: 87] <= in_ZeroWriteData[ 80: 87];
					if (in_ZeroWriteRegisterEnable[11])
						Reg21[ 88: 95] <= in_ZeroWriteData[ 88: 95];
					if (in_ZeroWriteRegisterEnable[12])
						Reg21[ 96:103] <= in_ZeroWriteData[ 96:103];
					if (in_ZeroWriteRegisterEnable[13])
						Reg21[104:111] <= in_ZeroWriteData[104:111];
					if (in_ZeroWriteRegisterEnable[14])
						Reg21[112:119] <= in_ZeroWriteData[112:119];
					if (in_ZeroWriteRegisterEnable[15])
						Reg21[120:127] <= in_ZeroWriteData[120:127];
				  end
      6'b010000 : Reg21 <= in_FirstWriteData;
      6'b001000 : Reg21 <= in_SecondWriteData;
      6'b000100 : Reg21 <= in_ThirdWriteData;
      6'b000010 : Reg21 <= in_FourthWriteData;
      6'b000001 : Reg21 <= in_FifthWriteData;
      default   : Reg21 <= Reg21;
    endcase
  end
  else
  begin
    Reg21 <= Reg21;
  end
end
//write Reg22
always @ ( posedge clk or negedge rst_n )
begin
  if( !rst_n )
  begin
    Reg22 <= 128'h0;
  end
  else if ( | Reg22WriteMask )
  begin
    case ( Reg22WriteMask )
      6'b100000 : begin
					if (in_ZeroWriteRegisterEnable[0])
						Reg22[  0:  7] <= in_ZeroWriteData[  0:  7];
					if (in_ZeroWriteRegisterEnable[1])
						Reg22[  8: 15] <= in_ZeroWriteData[  8: 15];
					if (in_ZeroWriteRegisterEnable[2])
						Reg22[ 16: 23] <= in_ZeroWriteData[ 16: 23];
					if (in_ZeroWriteRegisterEnable[3])
						Reg22[ 24: 31] <= in_ZeroWriteData[ 24: 31];
					if (in_ZeroWriteRegisterEnable[4])
						Reg22[ 32: 39] <= in_ZeroWriteData[ 32: 39];
					if (in_ZeroWriteRegisterEnable[5])
						Reg22[ 40: 47] <= in_ZeroWriteData[ 40: 47];
					if (in_ZeroWriteRegisterEnable[6])
						Reg22[ 48: 55] <= in_ZeroWriteData[ 48: 55];
					if (in_ZeroWriteRegisterEnable[7])
						Reg22[ 56: 63] <= in_ZeroWriteData[ 56: 63];
					if (in_ZeroWriteRegisterEnable[8])
						Reg22[ 64: 71] <= in_ZeroWriteData[ 64: 71];
					if (in_ZeroWriteRegisterEnable[9])
						Reg22[ 72: 79] <= in_ZeroWriteData[ 72: 79];
					if (in_ZeroWriteRegisterEnable[10])
						Reg22[ 80: 87] <= in_ZeroWriteData[ 80: 87];
					if (in_ZeroWriteRegisterEnable[11])
						Reg22[ 88: 95] <= in_ZeroWriteData[ 88: 95];
					if (in_ZeroWriteRegisterEnable[12])
						Reg22[ 96:103] <= in_ZeroWriteData[ 96:103];
					if (in_ZeroWriteRegisterEnable[13])
						Reg22[104:111] <= in_ZeroWriteData[104:111];
					if (in_ZeroWriteRegisterEnable[14])
						Reg22[112:119] <= in_ZeroWriteData[112:119];
					if (in_ZeroWriteRegisterEnable[15])
						Reg22[120:127] <= in_ZeroWriteData[120:127];
				  end
      6'b010000 : Reg22 <= in_FirstWriteData;
      6'b001000 : Reg22 <= in_SecondWriteData;
      6'b000100 : Reg22 <= in_ThirdWriteData;
      6'b000010 : Reg22 <= in_FourthWriteData;
      6'b000001 : Reg22 <= in_FifthWriteData;
      default   : Reg22 <= Reg22;
    endcase
  end
  else
  begin
    Reg22 <= Reg22;
  end
end
//write Reg23
always @ ( posedge clk or negedge rst_n )
begin
  if( !rst_n )
  begin
    Reg23 <= 128'h0;
  end
  else if ( | Reg23WriteMask )
  begin
    case ( Reg23WriteMask )
      6'b100000 : begin
					if (in_ZeroWriteRegisterEnable[0])
						Reg23[  0:  7] <= in_ZeroWriteData[  0:  7];
					if (in_ZeroWriteRegisterEnable[1])
						Reg23[  8: 15] <= in_ZeroWriteData[  8: 15];
					if (in_ZeroWriteRegisterEnable[2])
						Reg23[ 16: 23] <= in_ZeroWriteData[ 16: 23];
					if (in_ZeroWriteRegisterEnable[3])
						Reg23[ 24: 31] <= in_ZeroWriteData[ 24: 31];
					if (in_ZeroWriteRegisterEnable[4])
						Reg23[ 32: 39] <= in_ZeroWriteData[ 32: 39];
					if (in_ZeroWriteRegisterEnable[5])
						Reg23[ 40: 47] <= in_ZeroWriteData[ 40: 47];
					if (in_ZeroWriteRegisterEnable[6])
						Reg23[ 48: 55] <= in_ZeroWriteData[ 48: 55];
					if (in_ZeroWriteRegisterEnable[7])
						Reg23[ 56: 63] <= in_ZeroWriteData[ 56: 63];
					if (in_ZeroWriteRegisterEnable[8])
						Reg23[ 64: 71] <= in_ZeroWriteData[ 64: 71];
					if (in_ZeroWriteRegisterEnable[9])
						Reg23[ 72: 79] <= in_ZeroWriteData[ 72: 79];
					if (in_ZeroWriteRegisterEnable[10])
						Reg23[ 80: 87] <= in_ZeroWriteData[ 80: 87];
					if (in_ZeroWriteRegisterEnable[11])
						Reg23[ 88: 95] <= in_ZeroWriteData[ 88: 95];
					if (in_ZeroWriteRegisterEnable[12])
						Reg23[ 96:103] <= in_ZeroWriteData[ 96:103];
					if (in_ZeroWriteRegisterEnable[13])
						Reg23[104:111] <= in_ZeroWriteData[104:111];
					if (in_ZeroWriteRegisterEnable[14])
						Reg23[112:119] <= in_ZeroWriteData[112:119];
					if (in_ZeroWriteRegisterEnable[15])
						Reg23[120:127] <= in_ZeroWriteData[120:127];
				  end
      6'b010000 : Reg23 <= in_FirstWriteData;
      6'b001000 : Reg23 <= in_SecondWriteData;
      6'b000100 : Reg23 <= in_ThirdWriteData;
      6'b000010 : Reg23 <= in_FourthWriteData;
      6'b000001 : Reg23 <= in_FifthWriteData;
      default   : Reg23 <= Reg23;
    endcase
  end
  else
  begin
    Reg23 <= Reg23;
  end
end
//write Reg24
always @ ( posedge clk or negedge rst_n )
begin
  if( !rst_n )
  begin
    Reg24 <= 128'h0;
  end
  else if ( | Reg24WriteMask )
  begin
    case ( Reg24WriteMask )
      6'b100000 : begin
					if (in_ZeroWriteRegisterEnable[0])
						Reg24[  0:  7] <= in_ZeroWriteData[  0:  7];
					if (in_ZeroWriteRegisterEnable[1])
						Reg24[  8: 15] <= in_ZeroWriteData[  8: 15];
					if (in_ZeroWriteRegisterEnable[2])
						Reg24[ 16: 23] <= in_ZeroWriteData[ 16: 23];
					if (in_ZeroWriteRegisterEnable[3])
						Reg24[ 24: 31] <= in_ZeroWriteData[ 24: 31];
					if (in_ZeroWriteRegisterEnable[4])
						Reg24[ 32: 39] <= in_ZeroWriteData[ 32: 39];
					if (in_ZeroWriteRegisterEnable[5])
						Reg24[ 40: 47] <= in_ZeroWriteData[ 40: 47];
					if (in_ZeroWriteRegisterEnable[6])
						Reg24[ 48: 55] <= in_ZeroWriteData[ 48: 55];
					if (in_ZeroWriteRegisterEnable[7])
						Reg24[ 56: 63] <= in_ZeroWriteData[ 56: 63];
					if (in_ZeroWriteRegisterEnable[8])
						Reg24[ 64: 71] <= in_ZeroWriteData[ 64: 71];
					if (in_ZeroWriteRegisterEnable[9])
						Reg24[ 72: 79] <= in_ZeroWriteData[ 72: 79];
					if (in_ZeroWriteRegisterEnable[10])
						Reg24[ 80: 87] <= in_ZeroWriteData[ 80: 87];
					if (in_ZeroWriteRegisterEnable[11])
						Reg24[ 88: 95] <= in_ZeroWriteData[ 88: 95];
					if (in_ZeroWriteRegisterEnable[12])
						Reg24[ 96:103] <= in_ZeroWriteData[ 96:103];
					if (in_ZeroWriteRegisterEnable[13])
						Reg24[104:111] <= in_ZeroWriteData[104:111];
					if (in_ZeroWriteRegisterEnable[14])
						Reg24[112:119] <= in_ZeroWriteData[112:119];
					if (in_ZeroWriteRegisterEnable[15])
						Reg24[120:127] <= in_ZeroWriteData[120:127];
				  end
      6'b010000 : Reg24 <= in_FirstWriteData;
      6'b001000 : Reg24 <= in_SecondWriteData;
      6'b000100 : Reg24 <= in_ThirdWriteData;
      6'b000010 : Reg24 <= in_FourthWriteData;
      6'b000001 : Reg24 <= in_FifthWriteData;
      default   : Reg24 <= Reg24;
    endcase
  end
  else
  begin
    Reg24 <= Reg24;
  end
end
//write Reg25
always @ ( posedge clk or negedge rst_n )
begin
  if( !rst_n )
  begin
    Reg25 <= 128'h0;
  end
  else if ( | Reg25WriteMask )
  begin
    case ( Reg25WriteMask )
      6'b100000 : begin
					if (in_ZeroWriteRegisterEnable[0])
						Reg25[  0:  7] <= in_ZeroWriteData[  0:  7];
					if (in_ZeroWriteRegisterEnable[1])
						Reg25[  8: 15] <= in_ZeroWriteData[  8: 15];
					if (in_ZeroWriteRegisterEnable[2])
						Reg25[ 16: 23] <= in_ZeroWriteData[ 16: 23];
					if (in_ZeroWriteRegisterEnable[3])
						Reg25[ 24: 31] <= in_ZeroWriteData[ 24: 31];
					if (in_ZeroWriteRegisterEnable[4])
						Reg25[ 32: 39] <= in_ZeroWriteData[ 32: 39];
					if (in_ZeroWriteRegisterEnable[5])
						Reg25[ 40: 47] <= in_ZeroWriteData[ 40: 47];
					if (in_ZeroWriteRegisterEnable[6])
						Reg25[ 48: 55] <= in_ZeroWriteData[ 48: 55];
					if (in_ZeroWriteRegisterEnable[7])
						Reg25[ 56: 63] <= in_ZeroWriteData[ 56: 63];
					if (in_ZeroWriteRegisterEnable[8])
						Reg25[ 64: 71] <= in_ZeroWriteData[ 64: 71];
					if (in_ZeroWriteRegisterEnable[9])
						Reg25[ 72: 79] <= in_ZeroWriteData[ 72: 79];
					if (in_ZeroWriteRegisterEnable[10])
						Reg25[ 80: 87] <= in_ZeroWriteData[ 80: 87];
					if (in_ZeroWriteRegisterEnable[11])
						Reg25[ 88: 95] <= in_ZeroWriteData[ 88: 95];
					if (in_ZeroWriteRegisterEnable[12])
						Reg25[ 96:103] <= in_ZeroWriteData[ 96:103];
					if (in_ZeroWriteRegisterEnable[13])
						Reg25[104:111] <= in_ZeroWriteData[104:111];
					if (in_ZeroWriteRegisterEnable[14])
						Reg25[112:119] <= in_ZeroWriteData[112:119];
					if (in_ZeroWriteRegisterEnable[15])
						Reg25[120:127] <= in_ZeroWriteData[120:127];
				  end
      6'b010000 : Reg25 <= in_FirstWriteData;
      6'b001000 : Reg25 <= in_SecondWriteData;
      6'b000100 : Reg25 <= in_ThirdWriteData;
      6'b000010 : Reg25 <= in_FourthWriteData;
      6'b000001 : Reg25 <= in_FifthWriteData;
      default   : Reg25 <= Reg25;
    endcase
  end
  else
  begin
    Reg25 <= Reg25;
  end
end
//write Reg26
always @ ( posedge clk or negedge rst_n )
begin
  if( !rst_n )
  begin
    Reg26 <= 128'h0;
  end
  else if ( | Reg26WriteMask )
  begin
    case ( Reg26WriteMask )
      6'b100000 : begin
					if (in_ZeroWriteRegisterEnable[0])
						Reg26[  0:  7] <= in_ZeroWriteData[  0:  7];
					if (in_ZeroWriteRegisterEnable[1])
						Reg26[  8: 15] <= in_ZeroWriteData[  8: 15];
					if (in_ZeroWriteRegisterEnable[2])
						Reg26[ 16: 23] <= in_ZeroWriteData[ 16: 23];
					if (in_ZeroWriteRegisterEnable[3])
						Reg26[ 24: 31] <= in_ZeroWriteData[ 24: 31];
					if (in_ZeroWriteRegisterEnable[4])
						Reg26[ 32: 39] <= in_ZeroWriteData[ 32: 39];
					if (in_ZeroWriteRegisterEnable[5])
						Reg26[ 40: 47] <= in_ZeroWriteData[ 40: 47];
					if (in_ZeroWriteRegisterEnable[6])
						Reg26[ 48: 55] <= in_ZeroWriteData[ 48: 55];
					if (in_ZeroWriteRegisterEnable[7])
						Reg26[ 56: 63] <= in_ZeroWriteData[ 56: 63];
					if (in_ZeroWriteRegisterEnable[8])
						Reg26[ 64: 71] <= in_ZeroWriteData[ 64: 71];
					if (in_ZeroWriteRegisterEnable[9])
						Reg26[ 72: 79] <= in_ZeroWriteData[ 72: 79];
					if (in_ZeroWriteRegisterEnable[10])
						Reg26[ 80: 87] <= in_ZeroWriteData[ 80: 87];
					if (in_ZeroWriteRegisterEnable[11])
						Reg26[ 88: 95] <= in_ZeroWriteData[ 88: 95];
					if (in_ZeroWriteRegisterEnable[12])
						Reg26[ 96:103] <= in_ZeroWriteData[ 96:103];
					if (in_ZeroWriteRegisterEnable[13])
						Reg26[104:111] <= in_ZeroWriteData[104:111];
					if (in_ZeroWriteRegisterEnable[14])
						Reg26[112:119] <= in_ZeroWriteData[112:119];
					if (in_ZeroWriteRegisterEnable[15])
						Reg26[120:127] <= in_ZeroWriteData[120:127];
				  end
      6'b010000 : Reg26 <= in_FirstWriteData;
      6'b001000 : Reg26 <= in_SecondWriteData;
      6'b000100 : Reg26 <= in_ThirdWriteData;
      6'b000010 : Reg26 <= in_FourthWriteData;
      6'b000001 : Reg26 <= in_FifthWriteData;
      default   : Reg26 <= Reg26;
    endcase
  end
  else
  begin
    Reg26 <= Reg26;
  end
end
//write Reg27
always @ ( posedge clk or negedge rst_n )
begin
  if( !rst_n )
  begin
    Reg27 <= 128'h0;
  end
  else if ( | Reg27WriteMask )
  begin
    case ( Reg27WriteMask )
      6'b100000 : begin
					if (in_ZeroWriteRegisterEnable[0])
						Reg27[  0:  7] <= in_ZeroWriteData[  0:  7];
					if (in_ZeroWriteRegisterEnable[1])
						Reg27[  8: 15] <= in_ZeroWriteData[  8: 15];
					if (in_ZeroWriteRegisterEnable[2])
						Reg27[ 16: 23] <= in_ZeroWriteData[ 16: 23];
					if (in_ZeroWriteRegisterEnable[3])
						Reg27[ 24: 31] <= in_ZeroWriteData[ 24: 31];
					if (in_ZeroWriteRegisterEnable[4])
						Reg27[ 32: 39] <= in_ZeroWriteData[ 32: 39];
					if (in_ZeroWriteRegisterEnable[5])
						Reg27[ 40: 47] <= in_ZeroWriteData[ 40: 47];
					if (in_ZeroWriteRegisterEnable[6])
						Reg27[ 48: 55] <= in_ZeroWriteData[ 48: 55];
					if (in_ZeroWriteRegisterEnable[7])
						Reg27[ 56: 63] <= in_ZeroWriteData[ 56: 63];
					if (in_ZeroWriteRegisterEnable[8])
						Reg27[ 64: 71] <= in_ZeroWriteData[ 64: 71];
					if (in_ZeroWriteRegisterEnable[9])
						Reg27[ 72: 79] <= in_ZeroWriteData[ 72: 79];
					if (in_ZeroWriteRegisterEnable[10])
						Reg27[ 80: 87] <= in_ZeroWriteData[ 80: 87];
					if (in_ZeroWriteRegisterEnable[11])
						Reg27[ 88: 95] <= in_ZeroWriteData[ 88: 95];
					if (in_ZeroWriteRegisterEnable[12])
						Reg27[ 96:103] <= in_ZeroWriteData[ 96:103];
					if (in_ZeroWriteRegisterEnable[13])
						Reg27[104:111] <= in_ZeroWriteData[104:111];
					if (in_ZeroWriteRegisterEnable[14])
						Reg27[112:119] <= in_ZeroWriteData[112:119];
					if (in_ZeroWriteRegisterEnable[15])
						Reg27[120:127] <= in_ZeroWriteData[120:127];
				  end
      6'b010000 : Reg27 <= in_FirstWriteData;
      6'b001000 : Reg27 <= in_SecondWriteData;
      6'b000100 : Reg27 <= in_ThirdWriteData;
      6'b000010 : Reg27 <= in_FourthWriteData;
      6'b000001 : Reg27 <= in_FifthWriteData;
      default   : Reg27 <= Reg27;
    endcase
  end
  else
  begin
    Reg27 <= Reg27;
  end
end
//write Reg28
always @ ( posedge clk or negedge rst_n )
begin
  if( !rst_n )
  begin
    Reg28 <= 128'h0;
  end
  else if ( | Reg28WriteMask )
  begin
    case ( Reg28WriteMask )
      6'b100000 : begin
					if (in_ZeroWriteRegisterEnable[0])
						Reg28[  0:  7] <= in_ZeroWriteData[  0:  7];
					if (in_ZeroWriteRegisterEnable[1])
						Reg28[  8: 15] <= in_ZeroWriteData[  8: 15];
					if (in_ZeroWriteRegisterEnable[2])
						Reg28[ 16: 23] <= in_ZeroWriteData[ 16: 23];
					if (in_ZeroWriteRegisterEnable[3])
						Reg28[ 24: 31] <= in_ZeroWriteData[ 24: 31];
					if (in_ZeroWriteRegisterEnable[4])
						Reg28[ 32: 39] <= in_ZeroWriteData[ 32: 39];
					if (in_ZeroWriteRegisterEnable[5])
						Reg28[ 40: 47] <= in_ZeroWriteData[ 40: 47];
					if (in_ZeroWriteRegisterEnable[6])
						Reg28[ 48: 55] <= in_ZeroWriteData[ 48: 55];
					if (in_ZeroWriteRegisterEnable[7])
						Reg28[ 56: 63] <= in_ZeroWriteData[ 56: 63];
					if (in_ZeroWriteRegisterEnable[8])
						Reg28[ 64: 71] <= in_ZeroWriteData[ 64: 71];
					if (in_ZeroWriteRegisterEnable[9])
						Reg28[ 72: 79] <= in_ZeroWriteData[ 72: 79];
					if (in_ZeroWriteRegisterEnable[10])
						Reg28[ 80: 87] <= in_ZeroWriteData[ 80: 87];
					if (in_ZeroWriteRegisterEnable[11])
						Reg28[ 88: 95] <= in_ZeroWriteData[ 88: 95];
					if (in_ZeroWriteRegisterEnable[12])
						Reg28[ 96:103] <= in_ZeroWriteData[ 96:103];
					if (in_ZeroWriteRegisterEnable[13])
						Reg28[104:111] <= in_ZeroWriteData[104:111];
					if (in_ZeroWriteRegisterEnable[14])
						Reg28[112:119] <= in_ZeroWriteData[112:119];
					if (in_ZeroWriteRegisterEnable[15])
						Reg28[120:127] <= in_ZeroWriteData[120:127];
				  end
      6'b010000 : Reg28 <= in_FirstWriteData;
      6'b001000 : Reg28 <= in_SecondWriteData;
      6'b000100 : Reg28 <= in_ThirdWriteData;
      6'b000010 : Reg28 <= in_FourthWriteData;
      6'b000001 : Reg28 <= in_FifthWriteData;
      default   : Reg28 <= Reg28;
    endcase
  end
  else
  begin
    Reg28 <= Reg28;
  end
end
//write Reg29
always @ ( posedge clk or negedge rst_n )
begin
  if( !rst_n )
  begin
    Reg29 <= 128'h0;
  end
  else if ( | Reg29WriteMask )
  begin
    case ( Reg29WriteMask )
      6'b100000 : begin
					if (in_ZeroWriteRegisterEnable[0])
						Reg29[  0:  7] <= in_ZeroWriteData[  0:  7];
					if (in_ZeroWriteRegisterEnable[1])
						Reg29[  8: 15] <= in_ZeroWriteData[  8: 15];
					if (in_ZeroWriteRegisterEnable[2])
						Reg29[ 16: 23] <= in_ZeroWriteData[ 16: 23];
					if (in_ZeroWriteRegisterEnable[3])
						Reg29[ 24: 31] <= in_ZeroWriteData[ 24: 31];
					if (in_ZeroWriteRegisterEnable[4])
						Reg29[ 32: 39] <= in_ZeroWriteData[ 32: 39];
					if (in_ZeroWriteRegisterEnable[5])
						Reg29[ 40: 47] <= in_ZeroWriteData[ 40: 47];
					if (in_ZeroWriteRegisterEnable[6])
						Reg29[ 48: 55] <= in_ZeroWriteData[ 48: 55];
					if (in_ZeroWriteRegisterEnable[7])
						Reg29[ 56: 63] <= in_ZeroWriteData[ 56: 63];
					if (in_ZeroWriteRegisterEnable[8])
						Reg29[ 64: 71] <= in_ZeroWriteData[ 64: 71];
					if (in_ZeroWriteRegisterEnable[9])
						Reg29[ 72: 79] <= in_ZeroWriteData[ 72: 79];
					if (in_ZeroWriteRegisterEnable[10])
						Reg29[ 80: 87] <= in_ZeroWriteData[ 80: 87];
					if (in_ZeroWriteRegisterEnable[11])
						Reg29[ 88: 95] <= in_ZeroWriteData[ 88: 95];
					if (in_ZeroWriteRegisterEnable[12])
						Reg29[ 96:103] <= in_ZeroWriteData[ 96:103];
					if (in_ZeroWriteRegisterEnable[13])
						Reg29[104:111] <= in_ZeroWriteData[104:111];
					if (in_ZeroWriteRegisterEnable[14])
						Reg29[112:119] <= in_ZeroWriteData[112:119];
					if (in_ZeroWriteRegisterEnable[15])
						Reg29[120:127] <= in_ZeroWriteData[120:127];
				  end
      6'b010000 : Reg29 <= in_FirstWriteData;
      6'b001000 : Reg29 <= in_SecondWriteData;
      6'b000100 : Reg29 <= in_ThirdWriteData;
      6'b000010 : Reg29 <= in_FourthWriteData;
      6'b000001 : Reg29 <= in_FifthWriteData;
      default   : Reg29 <= Reg29;
    endcase
  end
  else
  begin
    Reg29 <= Reg29;
  end
end
//write Reg30
always @ ( posedge clk or negedge rst_n )
begin
  if( !rst_n )
  begin
    Reg30 <= 128'h0;
  end
  else if ( | Reg30WriteMask )
  begin
    case ( Reg30WriteMask )
      6'b100000 : begin
					if (in_ZeroWriteRegisterEnable[0])
						Reg30[  0:  7] <= in_ZeroWriteData[  0:  7];
					if (in_ZeroWriteRegisterEnable[1])
						Reg30[  8: 15] <= in_ZeroWriteData[  8: 15];
					if (in_ZeroWriteRegisterEnable[2])
						Reg30[ 16: 23] <= in_ZeroWriteData[ 16: 23];
					if (in_ZeroWriteRegisterEnable[3])
						Reg30[ 24: 31] <= in_ZeroWriteData[ 24: 31];
					if (in_ZeroWriteRegisterEnable[4])
						Reg30[ 32: 39] <= in_ZeroWriteData[ 32: 39];
					if (in_ZeroWriteRegisterEnable[5])
						Reg30[ 40: 47] <= in_ZeroWriteData[ 40: 47];
					if (in_ZeroWriteRegisterEnable[6])
						Reg30[ 48: 55] <= in_ZeroWriteData[ 48: 55];
					if (in_ZeroWriteRegisterEnable[7])
						Reg30[ 56: 63] <= in_ZeroWriteData[ 56: 63];
					if (in_ZeroWriteRegisterEnable[8])
						Reg30[ 64: 71] <= in_ZeroWriteData[ 64: 71];
					if (in_ZeroWriteRegisterEnable[9])
						Reg30[ 72: 79] <= in_ZeroWriteData[ 72: 79];
					if (in_ZeroWriteRegisterEnable[10])
						Reg30[ 80: 87] <= in_ZeroWriteData[ 80: 87];
					if (in_ZeroWriteRegisterEnable[11])
						Reg30[ 88: 95] <= in_ZeroWriteData[ 88: 95];
					if (in_ZeroWriteRegisterEnable[12])
						Reg30[ 96:103] <= in_ZeroWriteData[ 96:103];
					if (in_ZeroWriteRegisterEnable[13])
						Reg30[104:111] <= in_ZeroWriteData[104:111];
					if (in_ZeroWriteRegisterEnable[14])
						Reg30[112:119] <= in_ZeroWriteData[112:119];
					if (in_ZeroWriteRegisterEnable[15])
						Reg30[120:127] <= in_ZeroWriteData[120:127];
				  end
      6'b010000 : Reg30 <= in_FirstWriteData;
      6'b001000 : Reg30 <= in_SecondWriteData;
      6'b000100 : Reg30 <= in_ThirdWriteData;
      6'b000010 : Reg30 <= in_FourthWriteData;
      6'b000001 : Reg30 <= in_FifthWriteData;
      default   : Reg30 <= Reg30;
    endcase
  end
  else
  begin
    Reg30 <= Reg30;
  end
end
//write Reg31
always @ ( posedge clk or negedge rst_n )
begin
  if( !rst_n )
  begin
    Reg31 <= 128'h0;
  end
  else if ( | Reg31WriteMask )
  begin
    case ( Reg31WriteMask )
      6'b100000 : begin
					if (in_ZeroWriteRegisterEnable[0])
						Reg31[  0:  7] <= in_ZeroWriteData[  0:  7];
					if (in_ZeroWriteRegisterEnable[1])
						Reg31[  8: 15] <= in_ZeroWriteData[  8: 15];
					if (in_ZeroWriteRegisterEnable[2])
						Reg31[ 16: 23] <= in_ZeroWriteData[ 16: 23];
					if (in_ZeroWriteRegisterEnable[3])
						Reg31[ 24: 31] <= in_ZeroWriteData[ 24: 31];
					if (in_ZeroWriteRegisterEnable[4])
						Reg31[ 32: 39] <= in_ZeroWriteData[ 32: 39];
					if (in_ZeroWriteRegisterEnable[5])
						Reg31[ 40: 47] <= in_ZeroWriteData[ 40: 47];
					if (in_ZeroWriteRegisterEnable[6])
						Reg31[ 48: 55] <= in_ZeroWriteData[ 48: 55];
					if (in_ZeroWriteRegisterEnable[7])
						Reg31[ 56: 63] <= in_ZeroWriteData[ 56: 63];
					if (in_ZeroWriteRegisterEnable[8])
						Reg31[ 64: 71] <= in_ZeroWriteData[ 64: 71];
					if (in_ZeroWriteRegisterEnable[9])
						Reg31[ 72: 79] <= in_ZeroWriteData[ 72: 79];
					if (in_ZeroWriteRegisterEnable[10])
						Reg31[ 80: 87] <= in_ZeroWriteData[ 80: 87];
					if (in_ZeroWriteRegisterEnable[11])
						Reg31[ 88: 95] <= in_ZeroWriteData[ 88: 95];
					if (in_ZeroWriteRegisterEnable[12])
						Reg31[ 96:103] <= in_ZeroWriteData[ 96:103];
					if (in_ZeroWriteRegisterEnable[13])
						Reg31[104:111] <= in_ZeroWriteData[104:111];
					if (in_ZeroWriteRegisterEnable[14])
						Reg31[112:119] <= in_ZeroWriteData[112:119];
					if (in_ZeroWriteRegisterEnable[15])
						Reg31[120:127] <= in_ZeroWriteData[120:127];
				  end
      6'b010000 : Reg31 <= in_FirstWriteData;
      6'b001000 : Reg31 <= in_SecondWriteData;
      6'b000100 : Reg31 <= in_ThirdWriteData;
      6'b000010 : Reg31 <= in_FourthWriteData;
      6'b000001 : Reg31 <= in_FifthWriteData;
      default   : Reg31 <= Reg31;
    endcase
  end
  else
  begin
    Reg31 <= Reg31;
  end
end

endmodule
